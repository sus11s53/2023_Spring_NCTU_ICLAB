//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
A9q3aFmf5loXotYmiXMC3C+10PIddaykKfgWksANzKCzg17vKIyZ9rQjyx7vTZ7T
yu/hSR/oK5E2SLhXpgPDjq2mJVybvZ+WgbpGQNExPTS/sdAHFizfA4PvfAeH7lNJ
Lzaot7WHl/ypHA8JbGcDYcZUSy/GJcm/mYXEzTpD6xCv/li/Brs6sSCOPyzFXnB/
N6OaUs/7wBFobk7NyX/8cDr3sg3c/lL85Lt8NBszHI7QMftTny3NcphC5KcKnCLt
HzrRSfUwT/VsFX5Pg0NXL9slkBgoC2wSe7f/0P83F8R/Oj/GeHbDoMghIbDKTYSm
L4YR6/FGRQCGIJTtbT7gLw==
//pragma protect end_key_block
//pragma protect digest_block
L7i7hcm6YR8Ldh7tbPn6/gcj8nA=
//pragma protect end_digest_block
//pragma protect data_block
xrpHZTOobauqW9eordyja7x+R5DBRddNmmbA44DJZJeP6lkUmnZRt99HsVWnrSil
CJn6zv/SvLEBEk+DQ6iYYeA7UVoB7MyrV0/xYjorcDyv9eYLbGcQ/Hr3n4PRb43R
Fd4aR3em0mycZb7eEvsFAI4DlwaB3yHxlnLigS0WPvCdx0m0dz6o26QWBfSWs0mI
QE9J6DNgNg2JW2vFAKAwCugjEi28gA5l7SsZUWAUthe2GCopN3GSqAbQRwdYUTLE
Z6lIP2E5n/5ShNmhjiT7uGKkR0EuWNv2EE0NjXIA7cDmCzhY0OaJYrzTRbklyQga
HORSXn7PNwNE5K6bQwmhulLxMQgZLSUTYlo56MYR9lwx9SKoeQthFI9M3HpVY+Pz
95cSJ2AYAt6UVmSyDqS47EagCHxsI7qpno+HDBGgTioVyxgXk5y+gYd7zIeyV0Bc
Cqsx0BAzNCFKJW3DcEXyf9OdACL57mMgG3HFE8pIrvm+oNXEfu21VlPnk78eA57l
dGlT4gSuIESJueGK6wXqDG953jsDO+3Ta3hESTZnZx4KIfU5MdjVAeimuxz91Hcs
i3Pu1huer/AMzeYGzp6wvfjYNQ5qIn3WPKyReZ/6hTVDoa85Pw29tCW+9KWlbeQX
QiCSfjuD4D6i56P0gosPwzk1umx+QS4a9AiaZ43johVnVtQGl37n31R9yCWZC+x1
r9ebRf3ZBGdGmy9fx1/Ako5AbdI0/d468v1KvFgAC0/jXRWPSqJkJTj1tHb0upc4
9l7vA20Ew/EwuhqWgGhY2vevRkiUja4t/JvfHPaF0oRd9pXyiMyg4dZMIOctQfmF
jXYleg4hPVWzlI2IvAdXHLiXljRk+oJ+uDPo7TbhBPh3lauCZhcvW23wlTCp/wy8
FKgnFTmUf+GcHDD4fmeS7Z0nnIL0VN/saZ5pgkB9V49KlViM/qUnsfcF4pRBrh8H
O33rWyQ+Pc31F1UZG8mrZBpu3Tzea80lk3yaeXeVpjzgxzpgsVzxIZ72fT8uCMUf
ahmwP8ki3hJQQ4dF2bKYzipciMrPwm8eCBpEScR1onYEO+ccQy88si5FbauJs/y/
xiq1xU+sEtaQ2Q82C5t5ovgA1J8ylTaeyVc/4zNGTJDTumJTzROzieC3En7DKkhU
7891A09GXmNsvgju26ZfXZYiaKJ+/IL7yOM0/cH8M10223VNqAp1qq8xKFPBId0s
vFyCCOQYjopvM05pTjKh6I/n9b9vPSDJseZYS37imjyZp57dMTwEBP0K5/p5Gc2a
bfrSa0H52fchJM5vez7fIi8eDL1ENXDvCboevi+r/Q9M7/vWJEnE9bJ3itHbWFap
HOiGvd49zYN5rmzjbCu0Om9JWKOf8AQtNzgzFNbHp6R+8rfaSqdfONO9x6ecr2un
GgNZZ1rJom6o0QoCND6v0dlL4EsoAAiwrXL+HEihay9bSr4V2PZZJA262xaeBkpW
XLpq40FGzJL2npNfttgzP8B5PjIGwevbdarfTT5WdR1zlrL0qvmuJUdE4YObLLsp
EoLIRuZ+St4jNLy/oinOGTx5w0r+pthNWY6qOyq3rI+VGGBCLi3rFvkslScfCjVS
FZPR7wB+I4/6e3EG2KPULp0EgGH+r1I0DBTGdlhF+6LcHfRZlt7nY2DD43haSNTp
3mEBPMbPvF/i/dzUnnTM1q34ALejzBH+1ZyjYYk0zpX+PeuhR1aoF65SgBxxPFHc
/JadOE1voNphhPMHURZBon9wZqXuy9YvCD6hAJjXOZaizaWakNUxwdX1NfNbhmmi
n6XpRvTwiZsbeocUGvJqVlv5IAxN77Rg/CZJkWcZumvSs1itGSYCD516JImt1RJm
d/U3VeEdETUZNvFK+KqyVQHG5vV4rydI27wBEc+xVOSuZaRdoQ+B4lbyDCo168oJ
KiLEkMbUR4blKSOhq4yI658RtYPHAWipJxrFfJWQIlFgKu1zfOxG4AJ2PzxVGs4S
rPFpx9mgOwv9U6pgwdNkMr7Yy07U6fWY75cn+qqclJSvLl+d0ZO6JGhRCwuphMrm
K7CayLR918v321t0Q3uVJ9b5+dimDwyxxi++o61QMsmPuNzJ44gelex2WVnTZWdu
TM22KHCh0tSF31kaSWa9HeHiKU67NM2H1edCxZwqXLlIvrxtjyhjahO86WF3ukFd
8XUri8wdcbsb7dnUJNTJfynfbD79cra8rGEaVt4nVi2mOBUvT5CXGFzco1e3OgrK
MRajqRhsZ2oQxTZnYvsUCS7+IS5ET9PjgbPk0C8rE18o++/KNuGsW0zKzwoQG8GN
pHeFF9Ps6Ga18iDhzd6lnlEXlu384QJ12sCzEJ9jwZHNmmHgjYXK7fyNSQBpINiR
i7AELpAsB/tPqmWncVT5ZD9op1Fqu0lDfp23SM8tsGAJlj9cKadSIUdABXPmQaYk
mfiHZYSOcGUCBbnqcz/N18N/G82XbFcoo796sQQbkyZkMTQ981yoD1M65IwqgXWQ
vQwNvEaDq2XeyLBSXnMF4fYRC9wMehI5AkFl0zXcDkFSBSrn2X/cezuMBN14a00c
n/Jb+ARh8Oc55TvJp9inIRTKUG0bo5nLpZajKQkq0Qgkya98BNKUl/9MzRMJ2tU6
xPvBcBX6VPdOfFFL7EycLlu+XdQ9F2AhdjTcGn+hBqwb1530UA56fCKAXo9iF/2q
Y0lnWn+Skltkxy5JxVMmQn0kH204RByqcIaLq5GmlxPns2FXSXa3Mb4oud6hHi0s
KEmvJk98kIWRcujP3sOSeIxnMVE7vmD7Xwrb2Lzexz3fyWmwmx8StaCzqOqqr9zP
AmeGWVsXvEZ6AZ/JyeFSp6YbNdufAe/7NSyp9rFxHEEcr3PDkOZ0saaJzLw4utWA
LWf3ikK08sb8DnqD+JmUxyve+1IFxKw7yO0yt/tS+DhxKLxs/KbpgS21DgMxGur0
hfFBX/oo8Zqx9taOjBGHkO58enY/0tzyRnmVIsdMoQwlaMqnVNUTV5yKbvZyCZPt
f51MSDZmX4HSDKmNimbc6HOEtp6yHipG5CnVjd4WOTV5E8/4UY0QW69LI5DfRJ6B
coYQt89b9fxMfB5244StzTsdC0yAiupmykNHSDqB6OQVjeY8nEwZSXzLdoyuwN2A
0E+CeKRicZhnqCkdC3pD8iJvY16G+u/FtqjAubJZs0gvR9fbzhbdgHRfBcPq9tX6
+VptaUSnnrzmzNabJAQIME220kdemwZyiE74cwA+ImV+raMya1cfsRaUjjloswlo
uAw6EGWWkYLvSARZCEY7iZf7Mqe1tBT864yEFcLObSr02NUHDKsM2rV7KE8IpThT
gBOLilqDoLk5T5eVbzz+XtQiXQe05T+rmDd7R/hjW04F0wY5MkBSYUn5kQrZnlYY
wiK4Xyo6ZYFXDxChBTB/kU0B4SLqWYUkvuyjN2X4mKXEvd8lM8TXC5GJ/jmox1vi
EtwU7wr9d54MffUBWTiZKSOszjVwwdjLGhl4EKEGigJzHHbL0fHlGOjcS51vE18i
UaW7hnN3h85hm1HZNc1yntAt9x5HpijmfInabu31S3vyfbh58hdjMM8L/0Xpq03m
J0P3ceeNr15mhRS59o7Vsq1cuAFYbAG1J2OnJwYJ1P9asvkYWZHR8q8fRPfdcjej
V7+GhgCy5b2zzyU+g9WWgzWJ4xfgC/bz+jgFpWlKzG/n4/Yre0X0Nbd8RNE2JrvD
rWLwehtbMz2PjlT0ii+80NI5sFOL/ZlotCOhW8vVsyyL56nDR4VAQhGt0l+a8Ilt
6/H8AfS2De8f51rH9EeZnCBNn2sLnMElEJ6ysgPe2tB+Bx19YoYwUF5xDB5raT5v
gmhxSFcwStdao/a4D4G8Fvq9l1EuBncUPt4lTXirbUWcfDfpyrqlHh5U2CulIFBY
NQGqOHuKPnDNf0RXWn6BE8WWgWam8ur4nDzNh9dp0pm9noq4hus03jpfzQrH6mjB
o3jtslWZasGzxE5J5nOyA3JCVl4ObwyDz3JPENyaqGx1YYKF/JEOpgYpRvnRW339
EG5ERuvuooXsWvG+oJLTQcF9VYaN1TwrDXg62skx7SdgD7TgO8mzmUs1koBgMVGU
a25jxuQDf+Xs2otkTj1bNz7ypzSXrvmhAQBdHJHu2dws4uurDmrZeB0Nr6d5Mzn4
JpfD5mnNz1PVp0g+9FMzABQYPX+bQU1MrHyWh+AI514Hpv9gLaMn9aIgnif9jmTX
ZLT4xkCKWChuAXv4fSn6HbQ8+Fv0WMh1jOtmi2qH6lQfkBnpvCcXzgofUHbMideg
0/QlXGGWx+ReEzJOQolnCiXMpS2pgMWvLPYkTuulbejvHQA/oOM5V/XgkxkMdMWE
erQVc8ajGFPk5tRZEYlmHj+GqeMToKUg5NTbNGdEvIWVmSWsg1olfMBGcIIFMYnD
fnxwH1vdiEdkIR6klziW1OCsbE4pbyWw1lPMNdYWkfwTQwf1eOoWnGbA4/88lWTP
DDC2qKIR/H7+AO/oaygqPF8LPKK5gAPK2Pfx/PJDADJGWdtZEDzz+e8gJDCJ1wth
O3lF3JRu8PU5XBIt2Vqu2/eI4y9BN+nU/hvqxG9BcsYkFbaHjX2Mdbcn2g4ZZ//B
yi+c5WKjg5q9YNC7qDogenHhuADuhcQCWjtoFf8b0DFQIsHENe0qr4JVhMvBucMh
3NC5F8/QSyVWCOng8PQ2N+G213crh3qioZIlwuNE3otgQ9ke6+RdOD0Juc45Sp0q
C+nOTDGQlyDn9h0BqSe4KUEuUmPUrH6cix3dXugSCCvVfB44sRqQeiKU38SqWXEJ
hQm6yK5WomHcj9ViqXflwe5pFuC1OivRs6bX7jrTmPzhqInV5rvn3yNzFgDSOFqi
byIqywUI0bN2oUpRI799O1LqtgG2w0wKHX/YnSu5BJCuhmLKiRuwCalgCks8OKYu
M0slo7BqE1YUcmVKosX2urYPF0OHIW1EbHZCqO7KXsIZ0HpsywSGTbq//2GcuBfv
4RyulDS7ReneUvNuhZM7J2HUbIbHxexRqZeowZibijDhNVrql13IonYC/HireDcf
BY2kQCosvI3OGiMdOxMadVyQPoUoGG9AZD56VY9IkvRN9joM1gSbu9nJR7BCRTf+
mvjkRJqdz/SaD0eFVqPA4E/ZhGOSvrfdcr6k8LDnxng1p2Cgn3mSiQ9zwu/9VoE2
2EpGaxgyUox2/EgYLx3N8Tuf6Dc1ebyLTYsVf4EzammhI0JVGFN3VqtTmAUL/CHn
hWW18Zwfoq1t2zT8YjAf5Fo/Pt4ka7DhPe++hvRBZdf6p877rGBJxv1QI8skWulS
UVXcBl2tT96Myueqe5+FUJy4ad+zmq4nYayXFGBg4LLFHJrWUgAQUHZH9SZkrVAw
7Jv/sjfojmJjcMLFWawIh4DU8TomzYtbFhmI1xb1jEgWbEpcYO9i8RQpZkBq2I8K
LWGZCL9BJAASjkSp2ic8VWpETfzpRqZ/kiIiEOpvNQRJxiqUHrojzmzfFnYQiDK9
/BmpXQmkPIC2R0Sl+WXF9dXNqKW3IIooqtiTbm9CB0WJ0NX+Uw6fTAtNKy9hz6nd
CqR858RzXqeV4XDTJD2bBqLB0p+X7wF64VBCfhYDYZjqFEAu6/dig+IWNI9DKh11
kUa2DDKIzBjGXoZZY0FvCMfQliL55KLZlggONLx50zaFC6o27mt1q2SQoqUZYELh
GG465xRT22KIxXFc6AcThn/CzOJ8GkthKxqGh0lYvnQbT+WHfff2D5uZ3rddKwGs
0594/cX8kMWvN9zfNGKGxM+CItFIWu/GRo6bjbwB40MYT4ScRnsjtqEzSGbLkrRT
RVxCVrWykEk9Qw+LXWUwYIZa1B+wIhtFZtr1NGtGl9jQYQUOX0SzsEcsm0oK5IwR
yE4PIrnqywR1fOCRaujuQ/VofaxT3gjsGXBWM91SUtLwMOsQqtgCj4mtndMoH2P8
N0oYs2llRYHDd2kSUP8EFxrwwJI2YUUpz3nILpEejzytHM7XxiUlyGkhCM5fcimt
JnIcXKEejqkgR+Cv9xMOpjOebzd6NXS8dRyNNdQPy34T/5SwThBmNAWz1M/X7i7a
1wiuEdMDkNbXE1stQYOScv/Ru2oSfh/t8lF8zDjr76OX/VoFSsQ7FlQ6e6HdvP04
rwc5I8r8xv51WVHYerhgu1tK4ikLR25f8lovQBGecdrf4g71hEphLh+18odxO8Yu
5BbNAXs49U1oHY1SkLYSCEjTGEG45isdKvEaKF/1R0+QZ74vUeblCV7oziX7yCdP
iy43CeswvJvuz0tgxZlCtKwPOeBVYhK2wcTcAqK2uOy2VVFwHWXcC23zTWzRaxHr
trtMgjyp6ZF6fm4iydJgIA5tnBnaxd68FXWROKX27UKsQEW9a26zFfvZMIqQrP7W
Wrgwl6f/x+RK5j+pYlsMqAYZ81QolqjwgBfD8DMuLDb1sFy2uU3RNrsFpttqUvfv
SNtdb5vLDmVOpFBF9aXiwUM561fUyZu1oRmOg0IgOUjVy0iZhxTMvQsOZ4Xv8OFI
2lHcs2ZvkC8zRTf/GToJUFaQLMXkB6ZajRhZ9AxfgASrp9ef6YSLubLc6VXbhd9p
5qSMxf+8uUDDfVDpXX5EJD9De48cickZfFfIhkedjnFdHGP2TFOrs6LnMBGOPoEl
+YMP30PjGIkwgryobV0oDG6SfC2l953JDAcFiYSmdBljFMH/zlbOlDgk1cRAxwsM
FjAaMiffJUSGihhwsSs/upnHbaNvXQ8kPJ2ZxPyXaxAOuS+07mcPm+vAxKIVaEAE
udEPwQaka6/M/fEvC/LdecEhLyLWfuMUH25O4EaqBwmz40T3UfkTlYvudi7MjPIK
wCmo2TI66xFUzVckfp7UUGvZYYrl65tiICKzv/NVCVJgQiqVk+teymlG9A4SveYT
vcysMQ5LDdNOxVKb0pgFnoO9oCoG6NtThh8FvC0zx6L8sGuOL9Eg7U4V5w5PCHP9
uw9Ud8FJAvL3lWjtPnZBZknofEjRrTgEinXgNmJ3KTfoTzDts5aWxbHBDdpH/9LC
zWeOmC7harBiEzF4CYDNAmGW8bPSDaSfY0V7gxFqtZ7XuFF5iTsdn3FuErdGM2EE
/vAa4gYN5+SL254zHUW/JGSPIXxwTrFfk2IOg01F6PFops1iP/gkW7SbN5SHaAM0
QzT999Xq3Wy14ffDZn3sEpSwY5jgOhr+N9kH7SmTHzokXL30f+7vulHmLqP940D/
TjSvqSmVa4ZyUx3WqP5Wp2Liryby2OkUUmHRcvIp98mvF89W532QCK8G3hHqcGst
PDgYyO9bQG6aMYiHZYYBsJ3AozGA0/2J33zfAG+KvvTYtsdPNpWVqmVYEPtyN7CA
lQWf3RA3ZU90g4dbPaoUJSP7MB8jaHAZaVLutWRxgodrkXI7g7zDLO5UIT57hJ40
imbW33vJv2LeKaQQpqByzrDLrYIilIjSFY0Gj64AJ8Fcj2rz1vuwaEQ4ocPHyDuv
AeQgxrVq3nurLN3R5xoqDMDZbBxZXEAeRD9T54rXwckeSaI/twrje0fVuECnrwEM
Vz2FqSQadV4bJXHNHIiWdjodXBR1EWGR9N7VbMxLWVlAPbclPtVKNO5+KxeRd7Je
vFRRaBHuivlOBYD8p9EwpZLBUsZU9ZAnBzOQUCW316OMkzHlFtK/27y/2nlXuqMo
NjE/bJzk6YrheN5ibIpsGyRawCl2MxIXNxUW0PX6ljya6Qi77peIXCZIUr+zQbOI
tMWW9Yo8oBVNUE+urSXlj2DcGKE1sfMfV/8xqHs+dzZz7gtHQthAxz6/beVUPXAi
+x2ht2/MFeBT01UQNuug3/Wi9Cvj1vvTtE9tfTFivZ90/STct3eYymcDu7Y0qLn0
D8B4ubSHBcHYvru19hUeXqC0I1DqDMnzh88ZxX675zg/Jyny0m9jJQO9TElxYxj9
CPraTI1YqNs6h+yhIEFHPYoYkM95KmWuEm8ix3hiSt+PA7hI3COSSEKKxMiu9lK+
YXprjYjyIKverzR1uUh/PZ5wq1LuEjXbgrBuY4eTS1+njs3IijVPuzVwz2afj4rC
1GSAhyszZlCJbvA88PWaBpJRIddOpG140+DvoTe03OanO2cMYtFNcGLPiMPGrnQU
cXOI19KGRbddNAp4NDEZoGE92liWF1KBUAI6TG609dGiJCLsgRPONUMTM5B8DHb1
aI3a/b2w/JDzR9cAhOoh8N+BIz37wvdfyeCejUKZsoN1wKPpOD0eeN2lZjUd24Ts
u9OuNZZMmiVLb6wFPbBBLctPbMdwBgsAz14flyGe4eNRl3Epu/G8VrMN1zJGhIXh
t3SyIZ9cOZ06sK0IBOT+o0SefzGz5trStQq4LTKrc2GFZKxWqLWlwzZvMn13LhD/
6nyqaAIQgxT7t/i6Td1UdWO9zDoFcflL5UI2CnYWFKUX3HmuzUjv+uqHzgq/K5Do
daOz7VMo1NXCRz8qTBcqjAPQrG1Epj0P2O7YXbFy+0H9kEPwpB3rlyDHUwWZdmgd
s7BGfLbDowHusy6GQVhMaDcaKeWLUxhHG+Y8wg/wVYF9hpxB2PksTmCj60i0c7ti
/GkbtJR/ewpGzJRrwlrhM9a6AOJZOBOxe2YY7Ad4INJSd3upC6OmudWgWR+xoRDV
nCsJZ2I2wzANlqe8BI4+CDtmsADih6rArDhzC0kHk8L/0WB1dy4kllVNQMUH3rpt
JNoNe5vQ2cqbf4tthID7bzWUVwaUVGqqBDAVqSZpDNZedaZ5ziia2oyiOXCZ+Hjs
nc+uEX0Ix3zbw8AXFRX6KH9aI5ei7dwtTGA/+ipBmpUJmOpgpD1RRBDtCD9CkLFe
HL76ei1ZZyeF8gC2HZGTAHd0n6Rdc0HSY29eCvLnzxQOP8hvKRHDQHDReP989OuF
gC7TDzYUUtltGDTPqkRhCERf8arpcfcqflakHYqFOlxKOeCf6eIRuijpSWc07vKN
nEZztcIuTW1ib0lkH0Pga61/Zu5Aq/D1SVE+p+FkMfGrg10LCo3aVvBjSb3d1FgX
g7xXLmj18inxNkNDiWTiEcgBA5rkEdibW6aNMbL4lAzCoXw/jNzgDIxBC1yveYRa
0Kk3S5e734Rqb81vzYwMX0evsgk3P6mAq5oJES/gRQvPrmCkNFaH9tKpKnBDnhOZ
K3yUhd38hkU8xst5uoLTj1nPE2R1wvbERyQ8HbMm50y8meZ903HlqxO4vBWjqk6i
SOYnIkn0dwIH3PkCURKagYobdOFe02FGeYlrlOCoxY++otd2Uk6g8lHPI9jZDuUn
T6pDo8ZNSVFCnh8dJXwCUL5WDFckm2OVpxrz/Wh7oMXI0WAp7HHoPSMMiwjCDKrs
vs5U7gqRXke/RoGB5J7DcQpGFZ1gQXH7xkLqHtimQDWKNvn8hT7SMU8iPVDVoHNE
N2FaORUytoAMbHANj8ayf04mRC24Sf5B10V4YDQWj+Nxi1Oe0utK/6+7cGvbAOnk
eI1dNuMkjxjy7oP+lzuFhl43lXZ7fnHtn3mTPM2XCIkauXOIGPmTiGX25irVuZeA
v8BtrvbOCyhZ68OD2PGP5vxMGSNmJahHN79AxCRXl+oHMECqT+d2QSb44ylLUw/y
5vA7I8pQm0Gcb8p7N2j6ZTh9rQuZhYVUSn3+m0KsgV9o0F8UXmO29YZn334NsVFu
8tZHntQyFXlNwZYfhoCmi2Ae/qMWtiBCbDQqRBoq4j70uhCKJ0X/Z+RAKM5ZL9kz
rXtwtAp+zcFdXMQio+nXcK4J0p4txEiC/DmI9jl+b86mUlCc8yX1UfHSVGxVbv8j
5PGWPh9t5THg/uWFAAIonnCHLk9T/6gX+3NI/NOVgsELotfNHH3p0UpSIsp9ngpB
fTnVJ5WI8y0Zdkh32zHQCoj3Qrvp6G9pCR4e9G4i/OymoTtm9k9wTgPuOMqzOfyH
g/zkselfaOyiwLYAxKZ5fX5mFpgORkSnlaTs8o/Y28IIQzE7nVTNdnsdm4/j6KVG
1XSxVX351JKj3mnJZY5rQVQuzRt0zjQCww72AEK0P+S92ftGCKaXH77ujoHm0WGe
ZpuFJ/Ky3XzLE7BFhLeHDzV7+mICXKFhUcOmxUX904kJz1BbRzF1aI5C2NLTVWCz
p8+CSAVRhwiwkk3R8vYZvAvF5sURBS9zooQ7ozWxzggV93dMXqS3vL+dDpRfr3Lq
Jo9enlGBUGM+5d05Cih8yLWxTQonWRakm1pYv155htWcXaHDJufcWE/ge4aVDMDN
kXys9kwOKZ5+u5asjLUXuEDthkpO8CyLISTwbcPni/s38viyILfEZAq7YTrI26Os
eohnV23lMHgAo6eDsdSSDj4aO0DPpZ2Zrn7dji/iuKBZ+p6DZPo0e3714n+ZM0AD
4scYfSQQs0y72xdUi4qJezGxwapR0rzOvdrc+rS6nAzhsWrI4ft+sH+dNjB/Q2HA
Kw2bEo5BiQ+eDVFWeELwddAc0bWeWelOCbAS9L0FR0c76Frykc+JvMW8RMJnWA5h
z8s/CpTs9ETYP7c6/gh+e7BAA6G0rPl043XyjWUsMIz8OQqHpoGjUSvaozhQUaD7
URfus6QO6T0EC0GPWo0kuJNkAhdg7X2TPfAboXJMffkte9/Qp2xoH5zvWubngloa
B2Gh1ROiqQuz5MgKalt2BICRu0Z0tEems2zw7OVt7ZajlHpPXOBlxnKpu5aC9ked
iZw9LvKCO91UvDKTkIpbpitMJ7Sl6FQxw3Mg6+9kmolzYDoh45rE0oiwWBoLPHDO
HBaqBG0X01U686tUCRmjs9K7WpLPSsQWYJ7kH6iTUEFQsJmJ5wzp1p0wHcnkdlro
xvKlRBFmS9nYUMSBuWPaFcJfDtiyGnIF954UONLb5pDsm14s2mHdULWmdlGQI4WU
hmR0c2wkmxqJeEBeZQsGEWcikp6m4J8bF5zKJwLYxkPpfb2+R263UQilHL1+QHTq
VLEX3U+mEFiKIFVOq27SXJIblvGx4219zRJtr4PB7whESKJahXAdvzMZtnkHPADR
6RuM84UycMUP9Gj3gX9TYyVU2NF/+t6YhrZ3iPhUeKHvzJplGA/J+7is45E+dGUT
BFDPhaj1Dq7C607YDnWQS9rr/FvPjmfWvIFljbowtig2sMkdmRL5VreVkW6+EKV6
LpOdobd1C3vH/QVQ6df7n05Bh/buIgs54wyZyKTp/N3x6VNnHS89Hfn8qkVv8UFf
FBA+1gCJQ3wV7m2F9f+JSRfhEhMW8A5RZlZ8P+R+tKFWpz7ewx5NLTFFeK/fWp7o
JkgD81wNjiAe8U7DX752W0DAHTSHSvYmuJLlQoe3DWrXcYFwfJbyLgiBS+6SRwor
kGdUoouU4MzNwb7i7jwtHS6/65sBMmQ7XImJniLnXC9m3d5SsAweVW/udi/K+2vp
kLlCqjR6Kf1p1FaaBm9n2aPHL35Xu9yU0PMZnu1sjxc4QLesuryMo0haFHDnbKRK
AhQMAAcApaW/rfT+4c0TEdmdrRhx6gcoZljlwT7RFg9E+0J86HVtSnlzX30QyNbe
gjHx8NyDlV2xiPcoBByrK/Wk0/pNWRID0nF2YWuz6GKSeMOndL6QZgWJT1io6LZj
/qtloQrnNpNbTlPHvCTdjoCxx0c+MJMQvmhvsbS6mJmCwSsThBnBrwvlbwqVqNN0
lAAitSS7rJA5kAVs4EulsmtzMsmlr8GKZ6xDoKR6WlH80BRPHH8KpfwWjBDs4bP6
XowfSS3lN9Z2y8hCkRzDXgBuIkKiWt4zqQetcqLfmhCObNIO5KH1TTStbtQXbzBE
5tZwYpyw7VsMty3i+U6qQziFYSv3z949qHP71taTfJFO8cKe9SeKVZjDXNtnJYyO
xzSbJi6mmQpj4vL52h7zg/li6nadbo+PdR4ySGjneZT5/0E+GtDuzNmV1QDjYR3E
BgLs/vet+y0Hm/ZvasLI4BD7tru9VD0JsO0lIhQS9g/YEkYBhGY/sHu8PQ57u02a
Ulay/s0i+ZzZUHZ8b5D+DLH0fdtUzQdaYPaaaIMqws9Ivj8Rbt/U1vQk6kRnkXs1
WgMDOTIBaNqVmt5XOU6LGhVYQAS9BhL2781VVLe7/VcQ+r8MeIZt3+n0KqlTYYGB
R/vlkQxVY45Tisu9AMSI1Ti7mI/aXZV+RhpptF4SxAbVKjMxRkHRokNl58uoDkLq
j+P/UcpqfBMYs8qGhSKCx7DakV72mejzDwVIF8DvMJYJfQnSK2i4E6QvA7imGLiT
wUWE8xbbrIWDjd/QPIF6rwc2TIrQOyqbZ/2U4twDYrBrhf5G/PTUAxxIoFvLViCE
bjbo7Od8xkMwWn84rOxP7lgIPIpl72Qhi4FwvlPcDfYU9RGqnPN05P23ZLMJpRNS
p1Qg/V4hVM46JPrizJ8E8abDO+czDVqtkBF28DQvvIpOxOE34rYGeV83PFC5T1o6
2AQIGz5Kiz1+zCyIEN3Mz8JMXd0by8EKfpZ+uOhNX/TzyTymHjFXuMl3ekW3Go99
b8FQ4x2puTvp4UyUEDdnvwwEhKFw1G4FLRi2x9S5rUZ5jSH6EQZX9pm7ETqdApAf
f4o89Wu/XV9vFwp4hzt1QD9QMr1Vx9REMQX8WsNJ6IvinlZm8dht5fnIsM21mX7l
186PbRpWqgfBoNDRQDDJD72Qi5QRML4HgicH6599l2yss+4hE4OHei4m9WCHuRuE
kEqtVW4S9TyhX8p6pjA1tTCN4ZzRX/KSOH3dN7HJHSVXCg4IQ3YX3m97iYGmwhA0
56dAT25VPjUDEgZoctze5xRPLWIqg/wht1uXHaQcLrzGBi+70T8xS7b7ApRn0gkI
8XiiiilTkBU62ygRGU1+WA65H/PV3GIL1gaKlqBkcOk1YqRRpLQIaA5dCqln6nBr
EqQFEkZ2pXCdwgy5HAynMykpMYeo+qDMeT4+SteWV1azmNEczNbmw7ESB1GQqS3e
ParfKdhhQ40QqzFsxw+5Ra2I0gjRP1vdh6ZHyZCcU9hHLGu5f5S7JQH3rjyCTcZS
/rqgOUkabpMkWov6RWW6iFfD7hLBy4thJFx7aP7O2zcWczfSDmpVJ+9TWDM+2CF9
kc6apF2XRd0g+9jEBqTVWoDtlDEh4rPSkAXTqYj1gWF9zvSATMTNKnkQSGqEywZz
mGJmkTI4H8xHRmpUDNCIcx9X6LAz5JhnCNA1qJHRAISPrQ2MMx+FoW4+kXL1uYgS
mqPskPPs+GHF2v95S8Jm8p13H1dFEs6vGGX9/XgG0DzWJv4brgQIWKa2KRpgE633
DVIyIehCoxQ6PbS4FZZj8SYRh/dOKk0CyQcIDhxLI1+z9m5lLCQ2G0kaS/QuoFQV
PZ7Mp0aaLOuFhvxtLRVo/P9Vqg+1zFXLWH4cPs3qJe7hVus33Ct9Q/IhWTsylvqr
jfqowfPErgPOKBeohLqnu+UCfXa+cw7U1CSQNT3MtEtF/+tz45P9ltMobCoglkKH
Amk5sM41rtEF6n3h7X6gZj/9+10tjhHz/ceJmyebC4VqA4xa5pcSb8hTwnyRauXq
WNY8YsYuE5buSiY8p+8lRb7LJPxmwT/048cfy7InSjvVyee2FlBTJKdb39WW7ueL
hO7ut4I1CxUwobukdbajPQf3RR+n+/z24jg1vaWE6wpl6dRHruFlZyHN7YEtTWZ9
REg0h9xYgLRNsh0Ou7SFc61SJMxF1wDIgbNyScKn6IPeK3uoL2Utk+cYXvzlug6m
CisLq0oXZxwTTR02/WGdXKN2LajmjlIA4LF5MAsupdb1Qrg9uAKyQgkFcEhlLl1v
Q7lHaXxU49k+SyYX89Xd7cHq/tdHSa9OxOTU4CHhBKha0KDkwm1OWG2zwbYZRJ7n
ssDH4nqxZH/dcfYDqxmBo2EEaaxP2kCNWBbaKnMWc6pOMqXZwP8vhi/qgRyYyo8o
5ypkGsBMLlgzf1tCYJNY/AeM2fqkxmB67I+K6LJSHfp96McHqBvDglFx6AF4bKbR
t3hnbwdE7rhoJ+XgHiUSatPreu34yiVxzdLN1BSypUa3LUcoMcsrkd98m2Top6IU
DO2+1wpCAMCg3Zt49sS9zt9N+TQphBBOG53Ek0UPrnocn169jyue+vNSJ9V+XQIw
KzANzk3gjnMwV5Ha58Ihgw0xoySIVADR42UmW+q9iOYEEqVcFIw+cne72UqPOKXu
Mzj/pz4/lj2SEH6j6u/NOcLO7kgUI5ID7Zr32/hCMvNBNmPm6gMtQbY+5SjcQhXN
RznMRlXm108B56UKCf6aj32eZw3nM7hST/R+vH0iYS/pjHRW04m4m6rURnaEawpS
vJaDTbiQ96f7fu/szlJ3X8b4sKeqYIXOFl202enKv1rFFkqAO+lJw2stQVNVt3pm
KRznC7AIzpXEVsgHcse1MPHF+TPugYnQCcAZXDevc08m2zmp0M1CJJ3wT0kaqRK3
lneF73CRYu7iIbvTYskmelJnV3Rc9fEyhiKSleZRKtuRFvi+J1AzYoBfgEsPJ3bX
Oim6npOBsC1DdUA4b0i2F+RRkFVT/c7OgmTStBLApmGptqnS0gOD08gm8ehpYPHh
7y9i/U/zgk1KTtst/ARF8D0lD36jH6LO0spktXgZuq3ysmtYHxga1GO3/EwP/fiC
M2ZjpCFqWVU3NaNZJcM3TA3LNB03uM1lnbuQV3MMotv18IYPfsIsewZcaATrT5vQ
XLmzCoDVqMO8JkGXitFnast1gaOAH3ewkmzY7qW6CHsxNVSMI9G8HEVl8WMc03qS
ewE8NBx1doGwuHtEgdjpgoJNq3dqem/VyjY85gWgbyYYqbKYqndmU+IUhjdoht43
GfAl7GWyn8/Moxav88DXw92Nem9I71QXXMezKRIj8GLpVB2EPBuxHk8mdBU6XLT4
qxsTNaTl8TJ7aYzspaIx1v98O/lEp+LhcTtDN7/kWyDU0fl3ezUOLUq6wS1oimC/
YDFMRTZ20tOHUzJQXkWiNxnFvOzLD7nLzN+ioQArJfAMmXGi6gaiJB7QOOSsb4gA
7n+UEBQ/KMlC9F/5bilkIXV1jm2xKCPkQ+f+iA3X+LnLFOuSg61peQGmKf0F5yoI
qD7aSKIrGEthSi8PbUzetyg9LJJaX3psdyaBkHJhHy7TowlndqEMyPDldrb9COs6
9pBGhPCKcCQA+mHefvgXav/UyOwFv7Jo4nY4KfxaUDRdTOa2tqsdu0ZRuo1swME4
1R0ymamKiyC2pwTyP06C0J20NIsqLE1F3pr2rnTGbr4/xLlGKaSrssBQ97vYukFB
hvLew5upWjB47nxwThggnHJZABWmQ2kjsVSXAJhOi7RcZj4u0qXPwMxfJXNuIBUA
jkEmAcm/dvVkqTbLW1d9/FEOQ+aQMQW8u6HLYmlQAVVWIkqneVvNJpbY6I2L9AV0
oL8OFwbDNMiEPgw0pxDDXP1nKqqsBXVQpxkjMR7w9yiZquxVzmh30PT+gmZXY4to
ur7KG7CoQal9KV8WMawZqQLe+bouV0veieRV6w2XIaGSHXbMNx0km3ao4E6waFi7
jy3aHbZ5IeMWoy0hDUXdgf1lZUKZedowoMmsWXtWPkdixTag2tk/lf6yUuY8GWQR
zQeroUnrPZzTMrO/JAHbWhWP+OZfDWaoJGPBrGGxBFJ3briSjcBKyVXOSjYNmGKz
+QDHQmn/Qzn15/xvWXKCGU+a3fHpVO1fzKx6TQG8P4aPJ5c2pGHn8dDRgRXoi4si
+MqYOB02MpHb3rvuxcBzCOU5x/kfyoF/324EI9s/e1CgeJIMMNzMA8Zq/FtFcHGA
pSt+L4X3LlboD3aSuKn5P/lVUago5rAOQMrpD3O8mxQWCOGCq+QfwJ+P4nyG5gzJ
9jM4GhyDkaIA7GOQXH1lEVXj81uogYN2+I/U8JxcmXl/8KT25bMoU+AXefDJvEo3
0s86j7TwDGSVU7YJhhkz+7G1+xDFLcJw8vQgMtoVaG99aAuHvmq0aymwERI87xKQ
+hmpoI9lqsAhGl9REJ8H71Hd5gJVG54YiNVjwGVnYERUTtqSdqASCANe8QUeDHRo
dmtfyUOB0ZWo8v5ZyiEWydfPidbAWhxD8A+9UUcYoRo960EfWtfa1Bp/REbi8qMT
+QILGi6evOpi610JjgeOgUJMzzn4n9sF9oL3gA6VAw1h2mpydigDuLqsGsF2QGpa
yOkZ5xFXRUBMWLv2je+tAGazDxhSVID894R2zuYXFjeCJn55FuWe0YUf8Mv2bFPP
vYnCIl9szrPN+L5FgO5Mi0T4giMqGIDiJIZbosuw9YmHY/rQcafBcm17s0HnBBPf
UCGW84SwzXCd30AXOUShKT0VzlfqQvaAyt1j+h4rwc+s6dLP7/2TAicoiM4PQ3OF
QJqshq5PNkvKRZo11Bp/9xoZ1lqQM1L0z2F1Uqex600Z+VVJgsY8bTH4524YQL2F
UqAuvr9TarKyP/ac5Sm5NpeEkkucviFOhJMwvFgASB24ptlQFB31chDS7vafyhHf
Rt42QYr+jo2rpocokNkaZOS02DitDdnt9lXmO2P03x2wh++ZJDVlYN5g9mZ4EjVd
SeM/R6CLRIs8ONUVNbjZcxiFE1aDCyEe1Kq83McGQ87SHDqbc+h/4D4GaULuZljw
lSHqe1WMCcuIS3V8WF2N3wHKi+eX68KPBlIur0UzFqTvu7d64iKkUJPUdCvz51Ua
UkAMXAtn07q/BGSQOfbzhqYZR4lXD8GENONQ8Y9LyNCyfssSnfpw86iGt5yRYaUn
G3/9W0QF5dwrPiwfKK4Qr2FItwjdPGIcI8ZEPMnIzWWbwfFOWsknXiGr8YaplyL4
DcTb941QhmxERCyoNUaAok0Znx9r3NCCNKBe6UN3KetREWU/req+GldhMkGaSgRS
zzWsEP6QbqRsUsdrayDhHVDPIvq9oO7ZfyMVdvra+y8bSNOClBepMZzEVNzB3Jhc
vJJ9TaqRUIAJIaaQ5w0OWWpsX1D3vm9r0ZGNiWHrPTCojqcQ3iHNkqo7tt7kRTut
02sb6KN9KE4zGLNLVKNCdT0U1ce8wuamTqF0syB6j6oBn9XhR8gts5GTk3GtSrEZ
3YKL/mmjJAtbyNfUJLCjNL37rT7A3VfSqOaxqX0qwen6u+vtQo/a8JeVNzBVab2V
K7f+hicMCzhCxuBouw13OxDhB2H3dkLeag+lGz1l2iJkMCf9ogTwbmaSgjDvSsLN
yDNIc9nsRbdhoTKtyfmNx1C2nQh0RODLxlRWz1ZPbIEphat0YZnQYsvPlcrkTgGq
t5k87EHVUCDWlMFYcr7ItGN/Ilyy+ENOVXn0h9w7lhXbvktzX2gSC8aD930UUHHr
jBuVkf+wLw2fdhfFn1Zcv7JRetVty6o8V8RDiDV6Wau2NKKXEFjrDZzV3H6eTmNG
HFB1C1m7E1FmVxiluruV9x5bB9HQBDKJpVpoKOjMMwG19SBrjjvMtNDoZav4Cl/L
KYzunACtwre9+4EwQxK3o0fnMMDdLt6Yu2wn+kmQi6WSpMgCuDR5gttPggAGoMgk
6GYMVqqS7JSdOecVajSGWu8UzjEI8KaP0HEIQ6G4+nguauof6DRNGRAp6LQWjXHo
3+7lxQsWddCLHzmPxjRy4Pz8WdRU9O6VddmAbcaZGfLl9UP2ESY6+zAfKisQmsGg
FXrvAtDx3biOo6aWfcGuqMDjgvMHEeU+zm6dwKLsh0fHYrEnAqYzw6EKewX2SGJU
/OZ9C0pXzFvMv6fobXsCkIyMDUUD1rOdJVzQPz6uXBQX/vd2BAqELao2+WsUgS9u
bysEeycUIRT1xrl+mIVNNcQW8wzXzLPR0PFnHPmVV/rvBo9PUtC8jjGK8AlyGxK8
mMjhyT7y/LCrUv6rW2SxOOngIz7Xou1QWzgS48w8mHbjhHpQ2V1JoGCu13/QbbaI
V4IPZDZDTMz4r3y4DS6yowJyaYr63sDKWVkYYW7ENCtX0iAGlvT521TLlm6HzrB8
CDXHH3fgUw2M2jpfnpD7khCDfakkdAn5oPLluljJe+XFINv/z7td89Q3dkWE3u9c
O0b4LVqp5SiM6qxMzlAnCOXb4PELcLI222FrgB2hLNOKRM1T8y2yjItNcw2HDJbs
2BrbGJJVMlhwOhRxrML0o1wHj8BTbiqG9w6ojRzrtQiYAaxx9javJSSbiOSTObnV
d0XAW0+b6JWIWs27XbFAzi2shv2ecpdqFSU3cpvfJkaZ0USXApT8puOzGGLgEfra
pPn8AhHYCIcEH8ubT+uEt/VcgsmNvWUD5YOekVOluywi5rm7fHl2n+ANzD8rq23R
fKXOSyVs1s0Vl6dthzD806twqxpQ+AhkF/cCoczmISzrMPV6vXGacfxICoNNMseC
4d8a3FjSMwPqFF2JdA24oBX9OJssoLkaZuU0iVYnu3slnUVEpDKxKvorv9rPZk/x
g8PneF/1/B/QNdNVSGW4Zzznqbe6HXAeP/mwkGgBK/q9n45fbO6443SD9Cl+90K3
MDlHoS8MMEgIv+BpSF/rqAxC0BncI+4tCMUj0QOmnmhYpr1Q9+L6R1VkzbbJljmE
haL2HZHjxi0lbEX8yoneke6ww6CkKJRHOkVL1Jprk+XtlOfqnz8RGkzf0p9CX0Je
nKTNGPaNsjngAd8X1cfiUWC14OwgrQJrTyVo+WuW8Y6kdAKR8u70Ngtw0otBzOTq
ziE5Lz7jJYNpJ3oDvRdvYXvsectpOdtbWpxhiOIhrqyilVDy2Z0knx1ual/wNLGy
LZKCZ2IKIieWyu8QTOT5xEGLHsF7oA26Ij2QRktr+cuBp/3bl7HlINEGL9sVFeKZ
pUyWeCNfCaHr9EHAbO/vSa56srMvmJ2wD2QC3L51rlnoUlTtKX51dCG2+SJZRaVO
SsX4JKP8txLge7TeeNtLGuhKGZvGqmkEb36X1kwtOkT9rZfhoC4azRGOAPJXaTeW
h1rWUz+aixSEbJDt2rjrCc7ltFTrtneJYSmNzkKYsMYmqLa8wcjuc9sFWw4Fgtwf
MTtWhIc9wmE9O7nKO0vwzbdPtpjVHJbB/Pnali0ehqTHNvNdbaP0jsb/opuddF1R
Ylw1SEeg6JvUajk9DuyAeZ9vDCPQ6JvXc1r4I8NAu/ZyJVg4jzuWg0PxNmhl5HQQ
1i4PqLNcFfOXq+dUmQXkjIRX91OArFQB9yXtjZL4b9M1OKGkDk4NTmI8YA+lduXH
GWqm5Qy13wFYXp1fi0MC9LIK3xu2KkFLZl8iYopWB5FVw8k5vd0VhQXL7PEXHVDM
Br4bpbaIDCdghkdcOah+oX+4BK+PhNl0TDxGDhzlC3QH5msU4XJfLePhohWhhTi4
IZMNTULmUtOlbanoD47f9O0yJSHTld6HyvxZnj1FAc1KPBcuX7BPETeGePP/tpQv
SNXlDPwLwcz2kGLp6ujOM8CJaCcCEP8nF5zoXDtrLhCl/u3A1IAnK7M8/N7GpziG
xuK5o6m0xjsWhL4kh4HrXiI/o9U/HzkAUv/SmpFaWnos7v3esLKZJYiPbQzJkAL5
yXXCow7xwKknYrX0BxRrKDc9+8pAAjKC38OGS0F9R9t0ZEaZ77oa3ilXU10otAZR
oEeV6tuhwtyaFlit+oXWE4/l+sbx7gBThf9tvljun6QSwgAfRDYp2faxTGE9bLLL
bAAo+7eVnze4QzWpU36P748I5t0Q0+D593OwaCMoAkKxb82hIARjAuzehT8ilGLl
3mmEMHUIetaW+N39muh1SH0DkYpdg18gZhfxgGIZm5ebeC+QZtQEdIC+HtFFTLVi
7Ehz6Q47+W7xbqJBGyyoWELNigQY8aIaQXr9ta3BckgtnRrYzzzS3rRyxvy42kZ3
ce0/cvfjdp3YNKX88pOpFdJioFIfiBJgJ4R7tv5y9cjlAzBdLt7U+uxkS/8WDLNh
y7AwwROY2sGH/oj3byE5nDiAjvNdu73YNz6kFWsuholSD9hC/AoboTXMhddHk7kv
t40WeD2Ud3fNDWKIiRX9Zsl6UkjWmXaL9bccDOgKUUvkHaYYQdHWZ9gef5n7wZ4l
6dJ5y0LnDz1Kwqz/Uomhw1POxDtdP2nR0igQmhMtv+y2/K4uleJ7IcGGpGPs3JNz
d+eknXwm7TethD8n2+eXXlXl0IDIsF6bw9C6tgWPqSGu7LP3b7+BgB2BAVBji5Gu
l2Q+Yuu5EPnWZbRA1sKg5M8rK6vs3nk5xtKCKywTxxfCxmqFfzq6enA3JjixT02i
6qLMM8+wU2KgGnyCBBMHb4PVvF44HCY6m1ID+pclCkJh/IffM6COznPXH3AcreSc
ayaKZVCDHczcvTgsW+KS/DZsW5XC+q/eUC9ILXg5YuVVQCQgZIOS+vQlVZUEKH4Y
y/Cex98YgN6zmOWyVjszVtbpOLKfVv3Zqd+XkT51z6rjxbZ7b4nz0r8yPCJK4eUM
tsyAsDskAtYVpdd6i0hWL16WPAj37saQkzc92EQ1AxBxi0X6HBlTJyOa9V/dU68m
zVgKMKgDoBHewTSu82c6sLpVinPHQSLowrKZMa5REhr3pKcV34Htk33HtoM/mJyz
fC5GthT9CQNQq7WhRQQlbRSbYfdJcdZL9mn7+DUXrm21E9nHMEbCrsh45R806z9w
WYeAEmWwM/UeaoDt73d7nG2z2XKFQvHJpI19Xc4g/3Wudf5PQHDLPmzfFR8p0gxa
y9hLD2sM5QoeUh45Eo4CVE/HiUGEnZ1uyzez0ETtOCzr33rzLKo/mjC4EmRQ51w3
41oFaRSEYvD/DxnQZivR3bqzNFPNoIqztwhk2iMkwbyofH13QZcj6kRAWhSlmYe+
yHuotff3cHc9+C+qSfwfl3qxLUNZmpzehfCNStiHTQDPpWaOGlhHIavXVyLJqyRm
ngxBJgEbbBtL9Kp4UdlNFsjmEOuZ8PjoLFFoyXrKhtL2znv/4nonCxhKEI7RZnP8
yLU5AIodE2a4Fgg+nxNBjMmwyqidM0MoWJ3OafSLdspHpIJgPjfBJHpcvJjAHwnC
3g6HSoglaOUyiFpbwYvWayYtWXHSSLTJXBi7kpJ5nyJQf0A3sWmsKSIu2bti81Fe
ymObYpB4en6LF1RWjEZsQmzoiCqUJZYDoXC4IRJJVzP9+o0C/H70Hz+8BdbFwwcO
VXsNhMBhklA//dArBKbT5FyTO8pw2ADGGRlcco58BaCH6UULZ1gypaFgkdSmKsD6
gwXVTq4YeMhOoNRSTjPv181/78P87uj871p6G+xPDfpxwFX4WpAjwM6xrzs9Tqtc
4Grf41Cwro/KI9gEdZSeIzb5XZBWIlMoZcxq1y0iPVdy7APjmHI4N1SlbuosW11+
c8a4lThx5mpBme7plBy+lbnoD8Xtn8cjQN70Jebo3OBxzqB70IHw4IwAsWbHxudw
u6Z1zShoAmnJa2wsxWuoIpEI9XLYrAytm14WlJNeOIxBrn9pDFF3Was0R75e9NQq
IL9ZoXMi8jmh4JpCWqSUs9C9qXgf0gAhIs1rAG3mOVuZhg6tz2hGJc2anmHos2tG
8mgiTj9xUAHKaP5DmjnxU3R6DKa7qotERr0T86JO7aBvxLjM+7bQCK44cGow+0/P
+YqQbn5axHxYctcM7Jn7k5Uzzi+3GaMZYKBitluSdnBOB8APy8r7vatQw+PRYSXi
DB5UCtKbgwhIweMIDmkcyAdhjg89bk3LxDROP5KRBytluE4mSlXj/pqn/7Aee1pk
bt64jN/tGWYhZqEBgZuR0pc1rt4QU/8lVPtmEWUBLzcaYSqloPqyhXf7m2F0UZhz
Wtd0NgeedgKJk/o3qL2oCYpMUnVSPL9LIsG9MR0Il7AJVNXu80Sqm9EdBssGv4S+
sk6+hQ9UkdWq7JpK7oHJ3dWeVtedad+2yG6TxuFsoW8MFF8qkpTRzwyF8o6pKjd7
8bKZqlgoxU4BR53nHsrLLoejIt3EFsf+KkjyObEYF39NUyjyYl/duvl6BOCSTP1S
hZ6pybT66LBL8lOTqsp773ugVKMq5+JzGY74NoKl4X2wcvTQ4LNGtVywYbr0D8K+
gA18srhS11Fg7tC/gDmqUHnPtUgYXxmIrgWuxwu2AJhD2AIf3gLtpYAeZWFuPpWW
0udqjmuH9lg4VDOCTE9Hcr6l3YasIYgG6qTDYADSOV/LJigexB5+QqjYkMwbGULp
cA94ns4kZJZ5klVihq25RmGDRwB8QICTVzFixccZ6nPXELjpRabGHPBd0K7c33n7
GxM4h/i9397smus6MERFaWyv3IhSe5x3f8Sslv5Oh5At5NGcULfQAxbjElScwL18
W3SkZ+f/bsTZUXBqDDWhpHJ7NFAiPIPypvw4IpEZyqeUczEJ37buWVGVaYdEG/Bg
HxkAOCAoZhci82Alh1VdTud+sJtYOtJNe9JLjST3polQ5NC34SpSitO8Y/SIk31Y
3Q9k8TKIKVqsHvPtt8Tpc5fXYbK2MUV7PO14zQB6/qj5DtvgVDmV2/0f17iSFE5p
ZNcIsd+uf+DoGEp6dJihJ7LAZ5/1E9C3G+XkHM8f3Ggko/nCgPSrUR+9cQr+VOGf
Tw9Sm3j4yPrj0lfQrq4ACOlHT8m5Qgh8O7NxUgTJ5+vceIVgv15qJsoZoIld4sp4
4+DfwapTlLwWOF02vi36aLsEztrGQzd20l+bIGlKiatP8r4QR6/VpZtCc/2AwN+F
1fk44lT13Hr+/G8F2N4vQD73/0TVeLvQx4phCwQFOkm/ajN4xzNcXSzVsRyhN2de
GxsrW/YX/30be3Pg+E8bOFxqmD/ZPM/MAf6YDWNnOa5vIcNjBL+I8pUJMTM9dQoG
3gC3VMsF7q4LDxE/JS8TYTPWLV+a9asj7OMfhWC481t5qePp/HIvnRp93vFf/Vj2
IlGAm/vxX2jYB4nhxNuT26vrhlUhRA7KlXFXWwFG+sUiYeUoQkiDdfFNQJNzQdXz
tV6Xts/P8ACn4yloeqIKgukq8hhiA5NZl6T0EzVqly4NW0MbJBRZRXKP/5/xjED0
7q8zwZrRKYu7WXp72yjbkbfMIhhlyFgKWIyUlLVD3z459Mym3e7x2jTGWHVNvZDd
6Q1wftwR/frFnqk6+svXilBHWRySkBxXyRM3Ebazf1muCagjbWtHK3GIZh1zS1po
z9KoR+I14YVB2am/GS4/A+K1NUbKecSwQbUKzOH5sPawkotoe3baapU41tigT4TQ
aFhIMPOyQHSqkhc6oXZO93G8YKdhvnKynOewBoE+1UVkPRi0zcuNfrh832rplfZc
/4/m3NIAxHXqpeJiaOFEvZARd8HD4s8ixYSgTGWCh1nQUSSBM66xu+6qbLaPxQ1m
TFUJLid4Qo13AvFLU0LuQHhBq9RtEgzpg7Rl7kQ8sRYarNm7nIv8oInpOh+q5e2k
jZ9ifMz/Mj95HzKYH60+lvZdiliFjQryErjwyjrzrE9w6Ik9Zzf8Sh0/3ywbyjyK
rLmHj9rFFLm8PKK6faWX57jQQxmDGJTGeI1I43pUJmkwxdyZfyVDo+WhHltMVbzT
owXaJ0MdabGrr0O1JkvTIILFzdZtSJrHGPjbqLrKfItKHKQtADMz1Qrn3MoPkc4m
aHoit5Kq8zmOnXlRAGs/JGT4rG/CFJjmRF/MZgjdF1egBSvRnJUUXM6g9vXSFgNq
ahpOY/kDg4w7n3P46uVbTdhw5vkEQQlm7inDWx6bJOLGRoXQOYWxXHRSFWpV7PQi
B7iIofj8Qn6GWTpPIcM5XJMcoa16Lhqcg42gUuPj8dFmYi8V4mLMAe31V8aghMPj
tgXVwg6C0oeczcSel68gkwWhfV3xl3AtlzsamhyCCIebx/bQuh9q+xBDfsXvQ1iE
xTLy0kqhJEw6rdnD1Dp9p8Y1M4onzxlDg3RjD9OY1FUF9Hiw47HWrNRER9xwaZE2
QwVvNvb+egkQPhTke8aZC6P+HCypajty/0mnCMv3QT9rDioOjQTYalURpwUhGDqr
1yTDtL4eIIGmdddTzAHWa6I4WHxUs6m4eg71XPi0W9Te3ljPBD7VpFRHNLq+haJE
E1G68ANT+zZ46GR+HH6EcOmbdk3ao3W0NmdxD3VYoD6+6XALQGOdQz8ErUQuDgHz
Jnl+bDXY9w3vixsn5Oz1kyMOGH4eir8G3raPtt77nIwwFYnKfjLmZ1KX8fYJEWop
BUzR0ZtwitEYF+uzT4sGm7lZy4VSsuWAv9BRNKmYeDNv/v39p0nBgmz1LYy1qBnF
s35a3f4VNJz83P9MDL+WRzgs6MjnUGi7/gCZtuGAqR3w+ViVlNGX9MoOPGQNvEhE
6w9prNJ2/UmLLE0Wtan6YzHk6q5eoUbNb2FLs03jPuOt1gLAiK52Gca8ybUh5OBH
5c6FjU4GY6wji2VPI3l+EqztEkjnHK9XSlmM7FnG6RT2+vAD2JgaZJNhscQz185a
6XcqlJILxIipID5ATWh85nHKUAz9m0Bv0KEFstoEPE3nZny11A3ovZkwpyADEXI5
nARTeho7sAoNDyZRbgoe8xCzlA8gSbhvE8sOQZww1RgnXSpYW0jk8qoEn+M9WXcq
lvCP1dHgFzH9cJzuiCEQXr6/deKK+gvyuYVnBhMVUF6pRm+nb20ifwoQ2+HgSyIO
WWbPFotXLgCn3xprcgAI7Q+syR85XcYt4Cejt0g7o9XTK9swJ+5BHfdEFI7NmKHV
U5ETt4ZhOZrVP3J9Cv43gkFSGmpC5WRE27WCZYvD7GyMMNst1DBnvyKE9mQrrhvy
jqzRBvFH/DiloJ3nIY5XYwH6ayLho8hc/0IFtzguwXm7WDzWPbjReqjvbQUanBNP
oJH+wqZ/CHDQlSpOUOmQX+ypWB6o+bBYfXroxwJDCW9J4pFm3UhTdbhpz4UGZLIl
J3OzSF1hYXQ8RMWnMLSdgmKebmDYL7M6V7/MB9XTI64r+iH6UwBIc+/lW4A1Hp/I
sW1R8AFgulNKSZclzlbTz6JLCINBlgUhgcz2azb1rzH/O8H4aHJdkInKXgHRO6az
G8Ksszz9L3A+zCFOtfxBEKKKCT+qzgeZK43e/+SPNa6/GaNmyfYb7sLE4uxmiC/r
0yHal1muuUFfT3YEBvNhxKawZ8qopCmzozUOg4Y3OKdt3I0boXMCBCs6VBboTL8s
YcmV3hFaFqSmygOCyz+YVTNPXRer1RueUcxXF0ZU6t8qTcZGKkjHV0DOYdbwTZzj
0H6kUgW6FlMqcRziGB5NXEQrDOfVKTIifOuKJQMQYf4fwgORqLnW5rLz85J4Ox+h
Ko3t8bsgcXyzS6v5TE1EyKePG1pEoJ0AKB9sw1xlEaXsh8551KdDKZ1CYFezAfgO
Ds4zNx0+ZGYd7vFpp9peRnfELY21ODEOAx3ekKu007Q1ovgwoxoYKAwgroXPmn4O
cn33TnH5ZIfT5NJDWzn0riA41Pf7TGsrFoN3d4Mq3OyR0YF1jfkzKMiYkwX2ewAt
OixCdLjpx+FnibWf35FNqyJ5pKieR1SPqmgrTV3ZpH1Dl1MlnJdTyjRWas3/ya7Q
5p+YSBY7B2JeF6S1abmW7/caOMQrvsBovvmPnZU35bkwCAtbh9jjRe4cz5BGIv35
jKE/SgSC+DT9UFMC16L63kFWE104y8rTVlXWwvjF7XffD9H2RxOwTsKwQAUkRqTD
dU8jICdlxIOMknyBNVF92UVCqa0I20JhJ51UbaGLOf2k1cn2I/BLMn/vY7Zrv2gJ
OtvYcVHwhOOXGuItBpYYcILecnpdSYtfsjaGuBduO+5eRQNjy3WbwlP47Kt3w5rV
k/kPgB1L8lGYIBW7gGlLFJlbEr0a+MqsAj4XlNg2eNyXvCPcnKhw2otXq9ZnsRMG
fRJKpyG8z2rVuORbhXR07JGtk0pjprbBCDUUG/SW3jzwOjlDpnoJIm2hkW32UJmQ
+/RYRFd54frI9fea7Xb8XIgqKWBNkt8WX5l8pHqvcjO20lmufmbH8HFj8YKCU8XV
1Jyl6TKhmQCtHg1bEHT97zdyZJIlpPE8iQEQvQWhk8KuoQ+pJdpXNbGy68jtqjpP
XWOsgyLFQqxELHGnZqtP8xUECA/hZ4vv+gUPO4HU88nPfbt9jkAIJaq4e6d6FMGG
OchcYh6mKVa/F6tSchU6KdGMWskx/5puNmC43di4nJFRZ/OhPqIvQ7IqPo/uoNiR
sLF17AF0ch9pOjt4LcjclklsUtp3FH96JulM2uoCzG1HLLA16LykMTd9tJAm/rVf
RGGvrhZ30Qrr1Uw20lMA9ZZvPf+5kZSujCXZg/C1/nJu8YXxNbyPRIIRgmu4GuvF
ridBwJBkQx/lTZKR5lx/Z2wIAAtEw6MDvpDiFKAufAXYRZQFxHPjPpxVvs1PWgj0
Bih5HTazxYomeKjpsS/kgLFfqQdxhqxqZKYR4ya9BKj8mnsj7W3loUPorXps0X3T
LcNZmxTxEY30uamgGT3DuuSu3LeDb48oCHPVqWwOQNLjnBZB/6pX/4HBijgGqY7s
++7nNzWt/pYXKDsY7JLi7TpdHcSE85If6zAnptD957W4XYEGCg2oI4xXNfi0kzoj
PIbY9mhN5mK1fmuugIAJdHsZ32rmKYIQhsMvZmqmPy7YPK5eyH+v/Le4H6IulsQE
mPS8DIU0Y9YS0Ik3AANToGgSTsXKEctqdG2Ma5M9qI3Cf4yMK9ZT9HehbEbW6vmc
yxr2eRbg7NS1zmKdTGiDybxDxAQ8OzyHA/RZ3i6F1DdF/JVUlqHgaecGvSwR9bBe
a2IS+nEL61HIhKfJPLKxmIC9g+cJ4HJON947cTDAN3weqhQIi1/ul9mYIKpUyFjo
3G378WcxCfWWFv/hFWq2/TVJ2sAqkEOZrXSxVZ8DAOPYo7ooHPheA0JBUX+3A6Rk
D/icHvSuDu8Yxv3GJLR/QGK1+vB4Vja7s5IvCsOb2PW7rVx+wohffrcVGSv+Oyqp
wvJe8kgKXEJVJLiHP3IIlYabVcp2V+74zKHbg14kLCJiHWZ+SzdW8/vcgQl4hM08
ZqZnNclZzqglklHeO36lPLey6Evq2V4GZffUTNqt3SIoKQ0dD/ucUDD2AYaaRunC
BFuDWxd6A7qAGG6gX4rlIRijDe2VVoW62ZJ8ElEVU11gPl/cXIGO5cuw0ruJgms1
C2bGlKWTgcoloir5IWID0884tn/8pVYxRZOqFlE1Pfl8oTJYeqAXNSIcmot8ijl6
ect0O2JAopusaluWmsTa8OA47fNHaQwnqeBKxzEDG5W6sds4n4ShTEz7VpVLa+ZY
XA99p1oNWJVMpthC2/bOKw6JDJTShZWpTBbs3I8f0ZJJLlZIC1CKq3X74BQB/Y9g
d9tAvVb/AgEsd4sTvK190WwIdQSRdzFh2iNrqRPb+mPXvUk8/uWBkOlrVv9KH4cX
g91xXvCRLFtTG/vDi2pa2dAXntQj9dpXtebwf/A9jasdoIebAFwrkrEIpD5OKvvZ
WuDMofHhEQ/3MicAYBDpzO1wB1TEWgiS8zXNbNmPWNCXJrT/Y0oazOB3ZhqXbU60
/LhDBNTwpF0avvJ3/1ewjvr2NrO9v48frw7hcWllGAPRV5nV+MxMl7kh/ux798ns
ygttkdOyIznrreAyY39RJO8M4fcJR/2i3mF26lag1nFmC7a78fZpbtPHEU+qlJBT
yyySNdHxRWExgG2rYwlI4RxL9sfodopigKnVMgzkoeKUtu5y4QEc3qYbmzcOVIe6
+x//zdDY6/W5PYVBQAe9kZho+y1BKC9ca83sfau/MlAVze5yfdX997Que94hoRxk
QVBr/EzS9PKYTo9dP5WklO4q73x7bj+gF3Tj87tFm7sAj/ssxSEtoWzZKaSEqEc+
xr5gpdCP0IARFoomlTBO3XgxeI8ZTsSU31InBDL3A1BubEdvML28y+MNPGrbrf1e
hOyT+TYgubU9CN1MwnxqUqTNI4X2i08jxG/0FH8shLnkcOiWw1RrxwVBGMnDH+tC
qCxX6wVaioLZ3vkc04sYv8WE6zvlyQISrJZvp5ttzBOZRYSE9B6GBWLHfEas8Gya
5mCBG1EeaWkCWEsYTskIEOiyyIPmJoAZAiDtjDVibSMltU4Py0rHd8KFl57nASf2
lrmVOm5hvR8lKoEz3aOt6yLV9NLYvGm3DFvyTuZid/RtWU99MJIx4eJAf4BI4jpM
j/GKsIJ/0U6vnJmFyIr+O2sTL8xp5gZOFCaRUUDhM9TRGy6qYz5q5/FZ9CEMhBtR
SdjMofynn+hbDo1uiCGwLDkUZUbDGIl/CjPFK87m+FDYtS8wTjRNH9b8f7z37G4C
zz6YuJZDDjxjD0vUAMBUYFSS4Dalavy9GQJnQEekWGUkxRNz23OXfex/fo9oQNOP
XaEmBa225s/jB4s3BZZKyh5Hs6tyf+sX3E/6McmVHbyy3BdH9+koezdiV7PXxurj
zV63qfRp+bcyRVdxZ4gPU8WSmusc1QhWrSzjCZn3HsEUEgAbvgM3i9Z3DCFci17Z
DYvgJDoOZNseP1IjBZ9wEXyXsXuau2zGvQSOZU+tcFv5I56dZIYudjZ5IIjBYN+H
/Ntt8pODDyB734/qR4NEbrXD+O3BZcjZTeKp+Wv1yrQHbXh70uFb54+6PkpRK6dc
U2xpn7HnTT5nQ39XSfkUyF8G/Q52rNimRAQcRFLP3NoiHD2zcGRcdbFGVnC5IArs
mMTReo6q6lE6dCxG4B6E8Xk3mpw/DEzhISmfrkz8Py2cXP0SXIzrTpcyZQ4Y9Okd
/NebEWClM7amVmyTBODUNddcIxeFfySTGqsU8TufHA4oIzyZ4BfMQh/GfFl39ptD
DJg4SF/f32mSet0S0lG4dABh5KszhIxAXo+2ZY6/ZQZVrG8+Hb9njfyNedHKAa9O
AHPKvrZp2iDhpQR8tWdAKoKxGTmpnHpaUUk0LObGsKbveydEXCnuvpESOapBO6kP
VCNnQGUdfwY/J1+31zS5PwhdYM8kCiFiHpOu42GdpCchNpFORmzQvlccAFUmSLY0
ecWuIFFgJc4Jl3F892Qk8S9L3odqCZUHCLk4+MZCjKm6tDMtnh3LKeCIqjdLtqmT
Mo68f7fSI/FlrF7Tj0eRZBs9k0QBUtfKmYdgZMgwv9yiQhldO8jR0lYdipDK7xIo
zg1rHpHzrEeLTll+pXKGhKlpxC+F02eA28K0qxuGdPqui9erI8TeFlJl6J05ZuUC
TLvpxNE+BZR4zotsjjOMYKetqn+Ro6LqVJKb25cBDsrNmm9h3BxegWVKoWRCtQMo
vgqD+W5Dzj4dqLBdx54nn5bbafaaZvNi+ram7rRuSehkCCe1me2ueMuXex1TAUPA
deQ1doHpgBYWcNT6/PM5d7SdYkz/TwdTDE0wY8fVMlRPvf4CjP7ABS4gZjHpNN9P
ENT3XnocBAKs8fN+NUNa+VrcV0aFs2vNPsueeLDmccD1LQtOj4O+9uiBydXiqLnq
o36S38xAr1kGdT3Y0us5mTXTVmGIy8SA0FjwCvIrS+ikFAkTDrxvVdf/sAMD5cuG
e9Cx49+DW8AgtrFbFhInh1SlqXDldP0ysYoW3GeHlPlL0fgF7AsxX052tV31zdeO
rh7Oo79TQEMmk/acpx4ZWOaEZyqHKv2SVzI/QHr7zmb0hT8YaZu1n3FRDW3WGs1S
6YDogxZcHNj7NNAuda3ZgdCpcwOWOvAfuw655QwSQi/X9fJGrHuGMev0qL2UTN6k
snURExrnUJm+DhKE3H3smZ0a6e2/WzW1uAP2kjDUr8uYLur4HHQYGOcZ48DgEarr
dMjegXl7elcqyiEHMiETu5DOdaZTqPJmZarBwQ7WZWN9VojSmDxdIBRPHrbxFk3l
HGOnmLmp8zSYFcpLvi9TAKwP7CjXy+vr8ft7deI+hJU94WAADUHi+obBLhT4Ho5C
P4bbJGZPdZJUsdu5OqJjwDwL+VFVvqAfc18J6oqP4685ucl+PZLwPWLmOwT5zFlF
kt2bLqFbAUEwEESqnbpKQ7KOm3NLcsvmJUjK5iFjS6Weji7u5hYCihNlDSPEBj7F
vTCM3g0164TFqsWSpdY4hnsJWnjvdRH3yNyR9h05t8p0+JitpOFcFc1M1JqnKl8S
C8exQRxt7naLS3fk1mT8xNZYzWqbpZgBdkgHCWRGceNyIky6sKpSS6oPEY35KGU5
secFKZVDi1LsV23TcBgs5lOi1BJTBcwSCxM/CpndFOyqF3E41nywE5I5ahBfqJFw
ZGsZuX7rem79AbYjWrO0+awam6RawKviXtOsmrxER0ccP2kBHKMjMYh3Z0BHIpYw
sgsgsRPU3uTHZayvnjxLLI0X7ehVvSTQ3sBfJnsQQHNU7vUfarjjoDj+XzdPBoNR
LyOu7HWIsKnMpK8C35VMxeluSi36WBaZIN1Nq9d23B/LBFzqPq4LHFDbiQ2MzJDp
bXgyceNM4YWn0EDJga4DRcBTz13e6L67FiVlyMgR5pSoD/O3Cqtfy6p8WWpYmt/z
Em1U2qYufnr0NdURJhuSVX5DVCgnlJuUJfTv3rHCCnSIoOe/R8QWmd4pVx98CxBo
n1ZvTPQMq3vVOEWGhWOF+7p5kLZ0J9dbPVYJavdMtYClaGuiqDLX4cUnM/kZcdmL
9WjTNy93XSbNkEle/1wLUfswze/Y89MkBtCF0ypOssj9tPQIiFAD8hPKz39WRrAY
ZRmRifcj/OJwisEcKabNaNXjVj9a2JsdWsvMRDj4CDMek37HqRB432R22vMboN6u
GzFLRqIOeTtbXaQJcDge/TIHIqykIAQ/inLoHJG5MOUo2v9MlSNyjAxGcA3JM85F
OBapUDhnmtG/XujynFHt2TYAXJzC0bVFoae47E3cGrMvezDAl22Elg1OUqBYgWiw
huzCJESBquphAA34b2PNWjOT01L3Rv+5notQ3qu01OFEgDJGn/VL1zUdDBVzT0Ro
UoZrXpiFxGALTDxKHar/53qHXcVsiP0xPTew9R0GVKsP7siGfO9rXMu+gMITyUIa
oZTCmMT9tvxMWmrNxxjmydL9VW4LKfGdo3tYLVmXk3mE+U/G3OvOJJ6AZVfiBeIc
p6QdSkQ7QAzACyozUH32UYwXtJincX2S8+CL4ilSRt+xjDWnZr+h3sB+MHXaO+Y6
sgc4AxkURrdfMa8tnb+VBvqD8VZLRgT0nraxpLrWL5nDcbc01Ysw4CO0Rn0NTDS0
WSGjLzJ4bBZevVAWghdOTkh5jkuGW5s+GIBOWg2a7X7z2nxzJeuoJedaVagozfaz
zLilE26v4CJfYRNSxYlpwJJw1XvdrAFwI1NSSPsyk3K4Fs04C8Fcb4medQ0fH03Y
NJedcpw7F4v7JZjjrkT0POSsFKfwzXjLhsiNmKV/VsGlfy8m1oQbQL2btbADb/DI
Bze9d3NSfb/s9hsU/ypwM6cu1tdX4TeHGLxgDyP1MUtsv/KDP3P+tMM98xCCZZjh
crFXEObyPEU7deysYPHrhqhCNHfhf0f3HRwKJ7pSEaX0u2J48JNhLjlh5D2BW2d3
XKmMoplP2cwQJfg4xsZ/j/TAIA0orlRYU0QhmST02ERdM/84Rm/1Bw1oVn9GqjB9
4t3PFZV0BhF1QlA3Ky4tLlzfTDnhNVwoPjI7gF0JgEyZTYeF43+VavgIOmzSq1PO
uLSczpjkydAyyWC9Cibn3skybojNDb2XV9Fir65YTq17jH34oxJPCseKNd0X04Ru
/NMTzx7bbQCTrykCRTc6pBvGyhiIepT1CCsIv0GGWrcDO7eEIcWpgTJoQtaAmLqI
2arxwCwwDS+N/i934/aRKET8o3Fb/3n80BE+M1VujP1yUQaW3f+jFITiq6JooSx9
ILsiItn9+ZOlkqVD0xnNwUAWSct2ulCybhYpAXoPAjPVujQLblwC49T1OLvKfp6F
+CkUyHopFdX5gIy6cHD1TPL84FmgUZMn1wQkqFHyq3mePKkIy2ijl/2tOY46l7LS
NUSlQH2AE86lFHmILrHOKuG27DQdECOjduKfC6z7V6aKIzz+NXIwywxmw4w19A1K
E91Yx3HC5r4VxIDFZUTBWIh/fPwxtTAvP1vUFDiI3AXGMVgs8earf6fBgVr3vRjS
uR1I0keFz/aSQ1DcrxP/bTF9R4iNEsSBWZbnjF2EwVLndzU4dNoHb4QJZfsqdZKb
I18tc4upKcE9jnGywVVq7TDufnCr3v1005SA2RpDhSc2gF49/bPR+kDv8qvwZtsq
crsl9y00ZfnVPTeMi9swSp8rwfilgvwVCzc5yuYkH4ISB26DV2GPnLO2I5FlMr+m
N40JVjHmNDzjMgG7/jlgzubcyzepjqzKJUs8x3cUjT/4LkVsEWboav8T8PrsQcty
ML97g1VwSMN8FtKWmhFwnIOJ2TFssoCbH2VnMW1bBwN5q/i/dxqUN7pXOq3XLC9a
USknVrrmHYzez+DbSSF/SrqJoCn/j6/BGxYdc3wfWirtyEfttr+WHAniA9jdQi06
kMMCkHM5KbnLztKxZfzBCWSxGyAhqS6OCoa3J7LpC01aG7QRh1BMB9uzVH7aQ0pT
yjf1eYwQWviOfM2fE8+gzTYMsPHPHjvXnUwz8flW6jJts+lSCkSMXezwpIBoPQ5Q
gq9BJ9+8vgalNf5eHltS6HxGrf56kY+FwGGfX9tIsY3ut1OFwak2dn+FY9cwhOXu
kBvJlaDC8uZRViVbf/9mTj78W/4N47KfmQCIVrb4VQI5COu9eje5xiN+rzasGFmA
Wm9hqUfxBEH+kqt+Q+DzA/ndUHyHhWw397VB1fjwQY9unYVW8tR/Nzaw0naWvAgT
JCvkZd5GETDDV9P5usGy6ElyViqNway6+WmGAR0Djks9T2oPFaUwJSlIn+C7wMnU
vL4khHy1GhITHYQPVP7hMLd6yK12Y/fOPT3E/Jfnbrca/sFi8qfpTXowXfBcOJUK
OWCkFouVhMTckDUgVI9w6Go2SiK20T6TxPgwEhdgObNp+Qk28ywlMxMtWcdNVBtp
JBkAr6UMatZ2JyuyUNyJXcWpssq9Pf3sA273jBOVmTQC0on5h0ntvaKlSlYYpRcp
cTPEX+YAiBQok8LTuqJ6GXL0soqPJ7BYt0TWBEb998QUPjZfitgdfS0tF+fSQtvI
s1Z2iG9A83xX8sEc0DY6Wg3PdWv2wqHotl9o0Fc94ncPgfEiJKIYqlU5feyltP3N
lOMOo5YLk9MzqC3iOSxxU1j9QUCMXkzdWrqjKVVMiycFUCD38K4bkMA73m73c3Fd
aczfef0mVDDYHLPA3MnRw6FQnAR2YSPOa4mY5s1OuVD040cQAY2TiCMP+X9wGbNo
0M7CiqfDCkFCUM5dqmkIFYkoC/ByBwE7s5rz5DHS4Ms/wy7rVEzdve5tRxUiyhSD
5B9s6t0QhDzxJdCUaGdRWMh63GFKkoHn/nTWi05ykvzD+YAkDzji6fDJZ8KF6rTI
hMDnh1WOG5gY6Zcy5ax5x9A1+OIGulc7pB5DvTHKe4Aszc6qkIvQHmAjbVj30ilP
r62+yTfFlYjdb+wUt1M+iWap7LcS31NfS4pY9KgFxDbjsFnf/QZxAdBrHk8Cl5S9
Tk6OzZdskvEIk15fHTCP3QzYSQjIrAYs+0M6fr2fUO+KMTc7do8yzGptDYEcLTSS
hIgfKF9wh9zLx7lpAR7vaGPq79BpcUH5fahRxgAhQazcJBlXd9mAGdZ7ZqtNKHnQ
4neB4i92tIUyZeAorz6o2CZcqOE/4It5FHemA3SQ9sJZE2VGdJfmBEaLB97RV+03
UZrHQ0i6pSxFlEmDEor9mE3+5FbV8PGO/Eux0VmDTcqciF6kGxot6nbMsyKPBGst
YKoMGkIb0idiS/icFD0sWUREy/aA2NwNCpAY9GLwjYBPRtZGhuB7t8q/ZoYHCfZ6
V8TTEpCRtbN2/vSQFL9Gce5c3zqNLESmXREFwY71QZbOD7kBUBBvVk2sgZI6CxDU
Tuoe2eXBaFKrtXqmwPfBEjSDgMViq71FBlBHNkMrGB2JHrgqC7Me4i33jhyvTTmv
lwIlxaxNAuq+bDBA0TSYIdvoYj0NXbxRXhaIKXFykG4OW90dTYn+7m+uxmrWpwOc
VGyKY1mbtnyYX6BLkZGAWpW/bNiwiV2rN4ChkXBa+krf3krbVZ9NM71ePasynkEY
HAHewGEq92oRa2GDkpZ28XlffuDngRlRbCQNb4XlewKGtQuzXIS1siEPwJtGuthv
jU/jkXwtkYPGQCUKI6XkHS6zXJsDiHFyJhEzFBqdt2XhjvpPrduYKIIzGLaXw53Y
9gfHA5I4JxX+6KVCCcSSQk3JcScCH1sVllCfA2uzLwZnBA/7v6vSrfK43yeMpVqy
lOBxwyyuWlFOjL5WedW+vzZu2tAAWHmYI1fU8MTX9gWPpmeu4gUvrs5yipgtHlY+
xqqd1bx3xTTwhffyjgGtHt5e8TfFY1pSHPvBlzyZKyEt40kVxzSoicCgQOPCqLM0
4C2Q0fKuvVHGb5kjk2JuigxW5okYS4P9L58SEaB8pNb3zsVQEa7O9kOCiVUNAobt
v7yj4sF0xkRvc3gmE+1Wb6Ln5TLxrClZEsrS+1ox77sBd63iuUv4Dma9oLNVlujt
jaXIbgVVim0nDBlVvS4bq6tqzsmSuz76+1y2Mw4loV/TeOpaZd1eb63BZpY94d7f
hdF1I7FtV8OH6D9vqkeTMReDxDOr6dbFdKqAwBggwASGK6H2pfQjb/MKN9zdEUQS
evcKWF6fB2oeGvq/Jaf4zijV6yYlb2AEidcqneFQT4krXf7N3CF8/D4/AGhWn5Qw
3ApPQ20wy9kNo3cZRHPF2E5mzd/rSaJcGeggqXwQIfo02nYymjOuMxzBzZrVOtkf
CJwRBF2nf1gZAb21hPKoBEv7UIy5EFwfLWF/oMMXuduqNo03dYuYpD0NNgNsRWHy
NyXxnGYRdog/s3ZSdVYTALzukZhBjj5vwFopyxy9Aaev+kMd2AX5uNeFcqQIAI2i
9XdHMs/eseIHER9tQkKvKttowZONf2imkJluCSrpdQ3B2IkKAgScgm3XzwoCCn6I
R94x+EaJOVpwi7cU0KmHCUBbqrCer2TPyhkv7zbkacNX53bVJn1zeZDIkmSJwHFg
4TpOh/k+f3xf+2dY7WCwpbDESZc4Zofm5ghsFG6pwPlv/GIrTEcUDk1Qc2c6IWWd
60QaGpARrJz+ohfJspDpEI/VNxQapYoKBYDnHYxhZzdsvJHuAbuk/jDEEHNi1znJ
TjnL3AqeicIDALfGIoWDDRese3aNd0VkUJH6kUGDtEF67Yw6xkRFj/Nt8MhkaKC2
voOdqAxdzOJhvTCslCMOT5eDEnXxKJ9Dhv/1ig/2m+AIiq2JY8LEgydKkIWR577f
c0Tp7XoogRuuFWeDJH91QydnjEd2l52eX8/KCuVIIJWZSV0MUWjvJWvhJ9HnzIPp
rIKyyEqGD5TNIYYyammO8+wWG43b9vTYA0BRwkzFTgJsaXVP0lC50qSifWZeO0wE
lhSqYT4KfmVfFaO35cZ1p8/tr6ZQGieAD3C28mKOyAwIVoxharwJp6EepugnuDiZ
1sRYy5M/fkWDg1QCKSitV2DD0gPmgbCVucP/5XC+m5m8GONuVCa2rOZsMmoAYBDk
GmGtENEknLxWAZqfgb+WBcIiGnrVAcynmmx99Z8Q/CPPZxMvzag3rokcHtqGvncA
I5mELY4szeP65fNY32w/HcTB6ISHc2/0ROzk4vqOxrqXWEq+f9nwu1wMzDiiGGUg
zOgQ34XBhtrJhdrBIivhUSvO/eM1R0I+ku5LJ9CvjSHpQesOFfs59xRc207jJYG7
v1K7O+Eb8El23osURIEBgDScNhE1tfjaJwbkm1F2uuL/F53/0i2wJl42V8sLOCXV
txv9Brg7QQ+EOpSCLRqTazZDG4Gt2Pu783CCspsFicFyxx2lUPuGbMH09Fxr1pn1
MxhvALxGitbFkIANwKdHluU6D5PB8Bh7V5jsfLBE1YMWTnY3t2McfX4LFxPJLV6g
S0HGjYAWVlBx3+zVGPLkIezRAidKCgttnotjCRWAeyCMBb++oFkOJNpRwBhQUVyL
LDREgE0jbOt/ckXjri+gmKXovA8m7581XTpxRbrbA1xuckgpFd/GdF5jUX0J5E2R
ruED5aBWrDi9AMfvhcv0260ANQdfIWwQHV6DEmNUgxKz8vK6MSbzc97pu+Y+zPdD
CGVuF8a7z8OUzAcuV4Gge2PkIX8aWoVOuRieW3i2Gm3CCEivvDjsPnQth6oWQb73
sIeqHrxsewXAUkPadUpjq+cOeC9Rzyl6/jVyWJtHQbHu4RTPSAAs5v1USQOo0oIo
W0NNtk52dohj0r0hV5CxYndVkmLv+szIhG2/gFeTp1JR26YF7WLpA5btzPICpaDU
jsLF1A7+Edp1jsqxCyKEoPO39+gzWFoOjAhJ3SKVWfUUum++mLCV6IArs8fEdSyT
1XovzGCfVuGT3P4saC0OvocnVr0sxv6EscW19kpugVJ1QPMtjFaBp7/mLeS+IKK5
63erTk9uMhueL+RcAxzZjWqvVfGrPm14Ogx3fm6eHT3STQhTTMNf97thdfxlFXSs
8XHFECX52ffVTOv+bkYMocyvF+iZ7nAIYb9SVEvwE/RtSP7CdKlTERbPhdL+Iyjd
tLcSlQssXjqAUy8DWK3WrCFQ0j1Q9nMIyYRztRFdNQn7sfOAbe2eY8xwxsGSjKgv
OKcWv3rqfkpJfk/LvGJ+gDDDUWWzFml7RG66aGIGrgNJsKY+1Kox9SFgg2qNwBD1
FKfPuodVEKHWoyChUHygMvzFG632WF4n3Lod95ZjBeVODcedTR/c8AutwYYYN46o
hcxupNsFMQ6w4NsISz9Onzymr7hRXUZI5O3dzsByaZJnJgmSaTEeBGDpPVA6Iadg
hqYDezYQJFIgbiRC+M935ZY2CfPErlEtftAUOyIF8VIAeCbHUWbkvLH9HZJpgKTU
dtb9t4iQTdpgNhGeH3ntF2cCVOZTmJfqtKM7g3gtGDNEpbv4FkFmcWH5+eHFxeMM
ArkFmKLR363AxUag7sOP/EdSvrt6bXykxtqjVRV4OCKwq9jSCaYRfNI+E+1Q42m8
KCEqOKgCSvj8unuqhTaeZS7haKctqegZZRzxIfbLCcfUw7i3iXXYMrspM3BdOirr
SlkWXV5juCr2R0BN9uX7jTxU3AdxLjBRy+Gc+dcx1i465yf1YaYv6WRVs4mPMT9J
6yu7ugoCPBwcoVNG4TFcJy1Fdes4r5b+ct2Q/b7CzGZJ4qIyT6y44Vi1xDcfyMOv
rBtHIF4e+KEqIwYTksEwc8/Tvc0Yrz9zm7QAWHt1YmPUMgHD/sqaDHXse+gltNxW
P4nVHbj9NQX/DEPBn7w5WsvJeAS0MgvTbcs0a0zBbiAYb+6H94vrheBiAq0ZG64X
9H9TYalyDmslA+kRPTnDbpqkvLuoftvhta9Qqnjmfz2CeLRu96l5lAuzZnwN0d9R
HLWtybAYnLqovnHnPBdpNeXU8WViZdKbzT1wdbDWfsuqmQRJxtRCrt+k4xNJlLsS
gXmHubBeVP6hI7cNr/TKHedQwMiGB7aR3wdwU0xnZHLRRnU3S6/NmcA1hQw+ir5h
K41Au3Utu5qBY7ZjaUQ1x2qJUyA2rFYEqvBv0vOEaxBdUaqQNDeSc35M5GqGPHX2
VhIo+rpMB5OEkVe7JiTFeFujvCIZZcCj7XnZgW7Zn77F+5eD4+qFd3vTDTi1DdxS
nZRmiSLuz0T6yaV4Ttg8ll1MxIgAOHXlyCPcygX60OB01a7962btRzRoi6Hhf5fG
ojiy28PLqoo3pz5TOxqzJmjtSNKYXHRri3lRlStmkot/Fl8SThQUY4yft4uHhUIa
Y7hv3aeMJ0IOTimI9hZ+7biqk/HWgfLmpJtZgN6pbu4uJxa+ERqRw29c9iNTT2Y9
8KoRnzinlEda22HD9tV5rrE3quSXtbEduyXO6lyMJ7PO5CWOuy1gZEj72ABPyz4a
41r9DhCH9xgVPB2uw4TJBRhDYKteh/sjhpO9yoGBLxeeAy8T4cpqc2eHOaGA8KfV
uTi8YRssm397jWG/3l4Q2izrWRaiJK7p2+Lu53ASg8d3HC8ZvAu0a+eZxJBXHqS4
eGP44r0Wb6ahcg15nfv7cexsBtmqLmXnWXAz98Y8OqsHRDpViApkegmcNwW69Ged
YUSiqATTFxeNVxrqvc4lhcQ5f8ORZFNxsSYFVR5za948puhw+9hlAQFiSANz67Mt
cJ5QIk2WIkSj49m+kKRjHqlv5FyuZ4iPQUfVx1QmLKWbLQPrQFvAPquStbrkw5p6
4sJts/jteKEDYdzbdXI+ZQ4okFD5ugS9fcO9lakBxVnk0HiF+uO4+Nagh30XYDsY
6FqCyI9GncyGIWhVC0NGDGecCppq5JGrRPI8qvfan70qyvgJqmGrXe7/9aecNTDn
dEnAmU6DB0lP2KfwuXjgbxOa3rPYAjJVCxCYVweqO6ZWKIAXAGhaU+u7KB6Ohtlf
lq1RLwbofQnaYa9wTQUs3SV6152cgBnxsqzRMQGzMgWeizg/v6bAXQrX7bvrhjwT
oJaQmK8IWHzRvfLyFM4UoW4AnFu/fr2KFg8w5QDyIE7HTQ8wTbcsqdffY09gAcTA
jtQkqIXrdvT3z28UFpVxxD5/dk/8NOgptrP01Rku0nYcKmTbARkicvaT0Pq33oLb
ms/npg97vJ57WjxcPsfgdZw+BvB7ye3jjBJRpbr7/PT36Zp+NhC+yD3k4Z+K7Muf
5iFlrTaEwcPlwCHno77EEN5h/c0+21f4iWooxbMSgFmszeJ2Ip7vlkeMJ23DKUYj
vxjGi5XFPwprsbqfwye64FgNaHq5a5CPjwESRtUeeaRNWwCKHfj3f98KMX91USYU
ECr09j9d8z6zR3VqugE2R9UpNteDbFENEKSQ7Lx+KG8BFzCyiXjuITiMV7vKg7jd
DTtoMg8ghG2YwZw80S70KPSXiDHGGnd51rp0knNnvc/nIBhOFXtXLE7Ds7JOnmWw
MKEIpC8AATuOeInew/G5Jf8dSIjZ04R1czOohpTr4MHj+dc0470mu/Z1X15vSwF0
NyqPvRvCr/ywzS0Lgr0gu/SnB5Fi8KxikKml5LeHz8bMTdW9Aas1wV6PiwKMyx2j
R5jRAClFSE3nh2T4bBC8jgYjlWgFJN278uCwpkGqJoHkMKSKaUUhseXdUSIdbA73
G4b0Kacxa2FQG5PXoCY7vjf30SC9dYnnYPa4i/V45a3ZSRkNeXz0Mo+vkdH775di
MTX/SDhYQDXcRM6sSSuchw6vsDKxye6GskOEiw065A8E8s0p/mYAsCGBLJVWEUhr
QmrfvTXAN5D9O8chepN5sZOaFTeo8SH03WgZyo6rsEiKwti6lMLX2hzxcxfspk/o
1FptlzrwaJ98SwWYWufWz64zJtwHep1prv8MvIDAvvYPh3jRQcCJZ9l8qIaGjjgY
StieKQwwMPTSjcTwR36qB2zChqT5TbXxuRTWW644nm8tutEXB/crwkCSgW0NmLS2
b3WkK+z1bI6Xmqx+eGuE3s7tOd6uybDjwEKfdHziEpdDkjBmzSptVWVJ1PPV7gkm
dP1Clo1WvWRKzYypDOyoXxSdXxDbCtSPmlJKQL1O9bxVp23IEgnArKB786qKvLQv
3yJ2TGfbWrMulCCvRQlDuTrVKacEJsk4XZCtOFHn2eJ/C/r+jkJtQanp0Z+jJfV8
b49I/CinZOUHU3WPjlngW/4ypM3zGqMS3TavTg0SHY38G8EQufreUOV6MLhdVFCB
Bitp0G+EGSbBg32qB3k1c1U4XFUFuVxECcwd9Ble4C+4E52bBaBaFRDbScYtD4UE
2CbAUl6fsHZYnbdYPalDoYWGmR8WfWHBSkrmZ/6npubH6G29CIzZ9SJ5p7uWXgt2
T/mimFUZ6PW8fgSzqK8uPbPdwlvd4LJAYYYsAtvUQkpn2Csyg94mnP2q7xhw8/F7
AQL/7Zemfgs6bz08CO7u7etkT9N5onrAp0E/EqYjOQM8siF2b70g1L2HhV8EFmIp
QV2cAKOWEeEtvoEAjBsPcYY0YYWlh5AS3LNNOHIdNdxbY7kle2vm5GNJBwEnc8yB
h+1BeutCp7wjntfKI+Jg1qYYYnJW6vy75BG7H5/VeUAjRhmvw1TXVo2B819x2ri7
zxk64a2nm9JzYoayFcrXCK+tmHqVJYOlJ6TFCfj6Itrd/JskALSbBgTHOsllqCeZ
i2Fr08m77xZSehZL4bPMiM6gdeglzQHhZH//JvyE0LwgxucUXjY2LBFS8S8w0hlQ
bYqjFqzAeaMFoqUWS34jPo3JzUDEmUDDZ0cxsnM/3iCgLmXNCrELm34tAsfIC0lR
JHc9IJy80i9Q/aF6pbGkriuyT4Q3GjQjXAB035NvBOnXgySjvWAo1CWZJpWjGSuh
wSvMMMpQs7o3Ch2No6n05aBA2s3fq6I21lIAhQDkFS1AkWmryKHFI6ZK914BlHoZ
wZdwR4K/DOvc7DarKNlcXkVQ5gFuXbTMg40acwLF9etkBxTlKR3AafsQ5vdIuGZ7
a969ZFrbXil5jwW6EyI6nQhEllWgG0ZnArCaWzP9VoT4i6T/aXk/OteR//d4A24C
k1O9nAXiXgUhsSpoii5JQ45nD0LX72EukpObuk7mOfvxFk7bSnT0RzjSiG6tLSXt
RN53ivTbqdvO0LgTn9yX/RadopZPtBo2Rw2EavMvnRCc2GW0hon4q4BfGX4u0EFj
7fz/v8zmjUCA2W9ynsGW1k3NgFEx36rwK1GznpwL4FS50kQueHT9J0Qf28lYWtLk
WlqS0uAbpHlc8gDkGXK6F9nidW4YpcvtzCaJoMmgUDIZv4Cc1660Iijkbo5KQ9AZ
QZEc7a5QOFlq7eKjFUlO8WZ6GvfrnIj+r9l3Nz4to4s9zxAgU9tiQY00bfqDAle6
XAc2zX9KqSO7L8J4EOFK506VzNrOlaHH9RF5qLq28dDA+v90exCUkWolCPqfkoof
4zk6G5VArW/V+zhIKlCTNhXglkqXzPlOIYc3m3a6jqFyrdm+CP8lkaJr636K9ktk
Z2jmeGr8zc7e8Hw9PWk1FCfrnlU5S4t/Mg6AE4CL1ovKOAZzcyxGNHrDM61Vknie
JQGNHZxq3zYPB/ajQEe40Zbf0Y7l+GTd/zTQNPAwgVrnoVSYtrxbUcpuqTd0oUvs
EXMTx49lzu+L7CxnOX5gYscwB6Rfm9tEBlrauM6VlWBU/KEWuEdQXo40u16h1jl2
e16UDEh1/C+fgNFJuvw5n0AogwwNqneOtWTRWBfd+GHsu4reG6vuhofxO9FYl39e
3hqj0par9f17gV4kwWaDSrTwpL0pv+sF+bT/6W2on1yJABiwLIJzaZUJYON6P7BR
wiLxpr6Nu82qGSOoQEV+1+xiS6CX8ljL/yhqKddi7fJL1+/VhPyavwWtaOaZDb3P
iaY2atqxK0ndQkmoshMzMwCyYLNMpV0FMlWWjdivx63ENfcvifjvD/xurimZE59n
a0oYbJgrO9cOZjPzVHQ4poHrwFkpU1WwQ2A6rw31ifg2ZGb55Lv51Ovm3E8j+mIQ
XQXu5jq57Z8GbSavktb0+RXxvralx3gL3hQRZTYch/9Qd5i5+HJzWbN/yC9i4Mz3
kPTtt6E6Y7p7awgLzBsRBEHlaVC195ouGK6llwl6TN8USjTkb8p2wkkg+kR4tTY1
SKZ9f6aAoPoGGf00hqCPI8ruOeUofl72G9V8B9nibO4jFxzwKHdqy84Hy2AlPpn6
SNh/4wcOcv7QhaxrhaFWefSHR0N06rpxWwFmIObmm/+EAA8vhs8jtVTNRBsEpzq3
KKVdcDNcu2seUy55VH1tdm0NXtSWz/9gRCmLV5Myl0SHq6NMHDKstTlDhnNgP8/n
ku7iu1aSU8uwdJOpW+gjEDk0/B8JhcJM/mdJPnlD++eMWf6YsiKf4zs/G3yo109O
dE5aOrMOwvTPi5uWjR77DQ5mERsRpqwMPkolltQXVlVszoepmVupFzYrxKRSqPcl
swbP+ys8QMOTGG/Fl6d3qeQTJ175ru3ZP9dqG4LQ9Z0Tq7cFbQdDUXacklQ+P6/a
c6vN6UubHG3pxsu62YTy06yqaxcYjKTjKpSnbErUTkdhlcxPRcBdOfrfgg1uEHsp
3wGrNp9Vqi2OjTE6hX88bvFeTIa6FoQ5qHolG1MuYzTlAijfbe/lZ08QG7hzAiij
vDDKCwo7JfQ/uz8g7n8mYsUwQNKjZaoL/eoQOorE9+eteBiEiRZMf3o941vQ6K2i
IdJgB8+dm2afbT3KeBuqgDxe8hRCuONUsWbd0cXvLaRam/i2lnE4uf3MqKstsWZk
f4z6DcRFQn9NydjM8MOR3Aw0ozb2GK9qbxiaf2A90zhmXAAKO0z1jcF9q0tJreyb
kY+BpPHoyTokU4TYnt7/oF16roACKPNii7c0sqOMJQpAfc3KiBxqHH9ZcVxncAmj
YE07nwGdH+Oru6o+Tnsxj05m2sgUPN1Vsu4Mpe5zvCgxE5psk9jKDOtdpayVDtJe
dV20TUniZJvbZcDjHVLhqL4Bmz/VVYDcGWB0oCVINz1grxIxr7wPsS6oPgG4X5X6
zzonzbUSJX8+8x/bwo+nWms+g/8+Fb3e4QHHySFjXQk+gHnmgAtumwkJ39ZxHizp
Z52SAJ5iJVD2Ah1QKA56sbbWWUfwNZla3UoGbRpgETpSYdk3/t6axphQmZ78dGPQ
WFF62voCpR/o2EiyYBQMKWoIQx2yCajdFQfhkkmkHOL3Ne56t96YRHP2YGj681Uz
NOeZcAn4WzxnZbas8tIOE7D5YEEQzP/ftZ9DAWqtHJZZPjdf+7vcSz5HNcnmLnR9
/aBU2djWqSeQYnZYaRKuh9iUhOCMrWrstdyqYkhRUNhAV9BwufKG/NH0sLQorlp1
zIPsVs8cu9dxeF4mIHgbxAywnY5R5mq3iOlqPlwofpRKVk6sYfnb1FGe8QHOd3kK
AO04INl9ZTt9ujBXyJIbInf4tsWDRD6Jd+3z8mcPYQsm/wtvEiayJ2WFk54lPqiL
qC3aRZdjE/4KCN0F/McJlK4Lo43vFpHG0/TWqNEcIhwWoPYkHS8sJJR5i1De09hu
ocTJdIQNDhcQGwTB9tEsEoZsCR1AVxmWwNpWOls7/Y+5r9Ledq0ft5UJ8zQfxAEJ
oPeMYX6M27xWNU02vLYHkHtLjDW6Tnto6qXAi4uTBoQJHOj+YfAu7eyN7Vjs5t1+
aH/ziglIr15AoG2RBKXk3oP0TW7syYLUVnf/Cu+V+IIVOogq7AdYLZ+w3m8yyUtd
ZWKu+DZCdNsi6VlakjhCzUBz0WpHKk+GOgSxHBwIL/8uey7+/vzluYVuxU+8ZP0n
sVGoh/lFCq3bSBQdNPxy4lX7Tfipis82lsNPRg4XgrCWLDoaw0p/u8BIURCNk6gR
3QKCG2QroK78V1usZDweBewOpEoakNqtSoso1JWOeLXQDiWThJTA5K7AmpFoGTix
lSgdbTpTO58B3qrvKAaUnRkF0xxkpLOb9a6/uI8PoOHe9zosioJV9p2UEvfjTVNo
X7FgaDGDCdyKdVs4kTPyjJuF8jzmstU9bku9v4UjTy1Is+6LS0F8Vr9bIhoA4Ips
of3HPNjfkDdpdULzi9BWm6LEjJifznPGKISUv6EFPW1M/XGfKulTfE8RDFCJFu2X
sVHe9Vf69xpRWfsWaU7vSdsYIH/2LvsZVmdpmOingCDuO/i6sUTK6uHx+PvGoObV
iaJXplHSH3I3ReMFubokb4qb65wGEVn9twf8T6J6ThB14b8RkBDzrvOikt4/Q2yi
p30TmwT6NoNNa1a1WuO+T5ocG1yO+T4sCGRNmr0soB+mJT1wDq3ka9ulAi3C6dUB
MmX19kKMqkDY2CHDh6ak6Tn5AJlPldc7hmAR/4zcVVejzhX3oWHQBOs0ssuTFe9Q
mGTszcxsaISCLin4eJDqabwz/AGMRuEqh6lm9t/utUUEyHnQYWjRNsqGUIK72bEY
ToQBl8FEUphszzLzwpfFlSTa0kGiHyDRqsJdqVKgEl19+iQqcQBYW5O4xymzp6YM
+42c1JL4BK+Mb/sou3N9ROpaPnrTh2mq32QUu5sGoP5INkBhPYY3DS1ZE+WNeQLY
iefCJUeeisJAn9755vRifCdPBpAVt7Tcr0KDsITejcRj/LeGMIwmUWRSgfrcYtUx
7xlvft3HRQFDb1U61atVAsrvce183jK34flKF1T5EQrjBn/amm+N9TIOUGPSh6OO
aZChKGEtZ1m7xgb/+o+l3ONgtkMZfmI+EIDoAXowyv/EA0SBi9fVOSKuG91WpL5f
Ssqwvz1XRBGqOl1KNWrt6RoiG7rAs8cPbW8ROkAxHrtRjKJgjqPJ6nkSFNxp+vVu
EUt03RlCDGFy0/aM+Vl6tV1g2T72qntSZs4hSu5tq70onKskvI+fv5Soq/v54wmT
Kq2P3iX99+dbf0LehBLiGN4QzokcXVCS4Yge/FiSlMKBDnMe0oQH9SU+xOSupjq8
HzPcVYDIWfmWNPn1Q3eNvUuB5Uy3pWzBsPhrP2iB6Q8tDn/wGL5Oq01OYr6UDECd
2Ea9tGRrgZTqpwKvnWHgHUxnrv3NKux9zf2YhoocVj9CPjJ9FjLZTLUM7PtrliDs
jXvqIJUIbzuL5zUNxTOoZc+veeMOQgV9qGf6jNM9rOFfe6Yn9i7ZQhyDyGEZnmTz
9WIR7DeJi7fsSweSnAf4nNWuUJXTw2msm8BU/kdgDm6Q2PtssiZfxCrE04nSOxRU
NSLibVbIDFhZkBqk5aT36S3xknoqSFyhZVxmYzRll4aj/7NXdAVggSjLtZlM49BT
6whpzV9gXxit/I5pNkVfOf2PyqkvkcdKCbQI31WA041hRefdccQhQSheoNfy53Tz
L1xQDK4jHtMJyHYhHvFzvx5MdaXpFe/GZ797Y67F2uY9q0Jr0VRHhUQ4T+w+ro7u
JRTN072guEWhuW65XjEfZLI1/ePLzESBnL14QzpjPqVt/GH2pFSxdyZCxPwzWlI4
wYHklB6PDYLSZIg0PT5PgHx1vF9QRvWb01RMblbMcKQiGwpmp9qxMavRvctf8T1o
ULhVqtjRNLNCIWHVpTwvFUeNxjGLuBW2Aoxl0bbhnFlUTy33UJ0NA7h4R1FXHWBk
e8mcd+oK/R3H9G7Mdt+x0SZFh7uzZAIL3tuaUAQe5EA45mbzCCcmUcmAF4qkE0DC
1A3YgFz2B2IuCe1MT0CF8Y9XqFt/bHgdo36cTHeUYw5sIajqkAU+VjXqRhKNc1Fi
mHaettqGh/2NNpmRLbD9DbZOwOpomEyTyNlL6R602Eutb+LZTeQsv1I6npFb6lht
F3wZ7+00g68KfnTQkNLesNy5nBW2P742hVTYEIsg1sgzqoxU45+xYgpoE1319Ha0
xOGv8Qv8a3u/Y7a4NEeI8bhmvKIKxIYwlG7AKvrftIECFbt5UyDWPWWkmtxbqVZu
ZQ/fZwPcJy7v5RuQCFza65U0i3dvFPJMZRepfo00LrsAAtSL17Moahz5l1+9Ik31
q3ZZhiM/y8b7DPSgP1LEpFQH30KSkzUORM55842O5lxTRD8T1fJOmG7SybyGsW2n
KB2rqScZxFb9E9Dx8SZuRjXqSBZ23souGKu0MJYd8IMWMf7DjJNhzKjGDnaCwun6
CYOURBhwnhmta850Xz037m5YL6AwOrSpN/NNKOhpVM+EqYC6nxmeuERFTs/Lhc1k
cPcxNveUImKt9Fg9Oc0HoBDENFbW4wy6741KQ5d7Jd5Bm220y2pqO6aWDl37ZcCe
Q6n5piIgB8tvVDA/z/sF688RYJuwRzf0shIBL5TvzSgiqWqzOkZn2T9xId8ogK+P
N8N4x0CSqnMipXyF5hExSadwZQIqDT4G7Khy4MQSx4z6O/peMildr97Ani5jrzRK
CkL/8Yyyaa7avfeTFcuyQMh8lgXP1hpnvFrvKsM2sUFapFovlHfqNf9pNYYC17kl
AofPCIBAmrtCFVmRTG8GEmRfSpMhZvcFdvOD4TPuZ+Z6O1qae7ohMQLxIDTyJ1uQ
qfUF2diDrmuUz5dQ0j4ivbOhm+3Iz1XAjOiNVzKox8ke0lf0H7DmXFwxAoGnuX8K
E0n08BTCoJZ94mQHKcX7RXuNptp3ifsG53bCcPvjPJ+aaja2V8w2PjxHe8baFJ1/
otfSI0U0E9ImZoKGlkmA+vVasrqoahiu4WUUzIHEuRljnx6FG0m5j/lo6zqQcGmv
McLWC+MPLn96RfjteGEizrvYKIdjvYZOIKq895NDfzV9uxJIBsYKhrBSDfO4v/m6
uJtSzFVL7Xq3XfvBhUFRopTT3g448zotHh8nVcPk2ugEySk5YDZo2ZCFIwQQFppL
nRIQLdW9nG2PQGCpbPd42ZDFRgnJXSQMWsu097FQqerPcvJrqRByu98mN0M13WrU
GAcvFMPmo2t53kpTUnJqPiU5/E2EnoV9CsmwSK164CzWtRIz3VEGmXC2TzOUksxs
K8zcgDcWFzA9h68XK94M0ezG+w6kbdMebGghCFMakmpoREHJdkeph/5RrBOvGs7a
FaZKyPwCbOpWi/LHKetfgGuuTnqpKGxbEM842/MNXoJ5y/ZILBVr35L441ZgM74T
ycpOkwJ95eWJirmoyCGeG1CJrUT56TgBW6XzBy7cUYIOKrZIBAgdPgP3xs04Ov8Q
Yksb3Q3h0y86rL5Ap54HdrDAM1O2MumpU8PTu64OBgbJxXCjb4wzBCmoyMZbO9QK
O2bzYcHFBK56o68jPYqc+tuUHuZ5AqLa5vtcH/1FdEhqiv9dlsloatwpIvw5nDFh
Gc22xmRFQ3WWnVyi4izV8KYaWqSWo8q+Q65B7JfccIRdpyPnnk7FbTWNxTd/Vi0J
4N53eUD4YHiv47YLIsybik5X9Adv4zw/KopqmSI04CUewRYl2GCC+qU8Zkzwwr4b
RsFScMmytLDRenZ4xBXNN2KsWYSpkSeeSnfzT7IggO5RT8iMH7UiYUlIeKnW3nAr
v1SuPeciOhocobcqCqvLCJcedCLY8DrNpIQZlh/W2EPZDKspGLBH7x9BM5fuOSKo
/jL1ajI7R3iWHOgRqehr1eNBAsm0Fc2QoASWMkT6J3R18Zmt5BkdkTOoWpFJS6ET
27BrsNWizGmTzY3ke9c+JhOOEEuZlyzZjIDubFv3Yv30+Yc9Z2qrTXbP7SSFrjbK
BH59mPBOr5knUMhd/te0c+NBsJ93Buo1MsXlqqm2UaIM1Xg4ag3knXGC5PC0SWRO
/+xSslQ5xO/v25qWmkW0uMk9BkAIWv0ANvBTHuGLzGQOoTZPZqWnbrPYI28/IAap
eaE2h674j2+GU1J2QbH3AHAvI+/IEV7rLRbzSibBpeT11BjTu0ASM3qIzJOM7K2g
+DjLaX+U26twod0/2lVcuxggxTijj1sScnnPORav9K/vPL3u0TN8IeB2AQUTeRoE
X13joE60FOqPCypRCEwMWL0dIf2q26GtgXrPC4YZqs+O02PIaivyvy7Isqpx+m1b
sRK8OfeyoHpEIkRJmJ0cTkpGA0x/wXOPdCyAC5YTdYwdzhqo6Kgr887Z8iDrzA7G
M9l7jBLFT8N60SiPfXnLJeH+TqkwAfepk+EaAROIAqMbUH3SkijCIh+BOH9Ti4R1
P/wg/scdofUWRs8tp+mLgaxne9H56XjdEz0Emflfpzrns2C6s5ux1JLfYajw86Dz
8nmh4VFf21GfDViGEZswzQf3D/uoO+EsWj0TRH0lojb50XJTAa45f00sHdwOdxMC
loDxMPpWcaxFngo1xnesxu8B8OOCGE+tE1bxbB9o/75QZnOhpq6hyLvxptN9+IHw
qFfccZxvFOSs+rdbLGfo9QeIUgkITi03UmZj8orzmcf6C+8J4FZP82Rp5T1e2xYP
GZgRadPlOGJLShjRzfo7xeFxDzWA0aim+o1R12YLq0k4UKiq3ajHR1WJYUcTvSZN
mMrcjqMEvyDi3dFK7YTa1i3ym4hwd/wkWzLBTfotapTP7mNkz/moUNXPSWuzzdo0
ZNBPnskegbgfpe15n3TBfn8GpZQH1aRYLi7UEsigCr4Uzmt53HO8jRpD6pABBEVu
/A4Ppd99iJo6M+u5v+gYkOGAk5//rY1P86AB4T+usKbwWVPVqTwthKeseUrq7y75
pjBn+tDB6fvg20w6Iw1oQBdHa5G4EM6c3JRdx1QsI/bypyX/9b/UKs/kjPXeJa8+
RqOhAriFaoSDRUmOmxK1647zUEC4USfuZjMkLpOjgJ4wQ98rJIQNBCHMjzYfdba/
ggvVfna//JitBA0tpefDN0T0qPxdAkzVPNrEXQ11W22XrbOeOmy8R9lTkOHyoNpL
FCyiw3hlJ30BUjKNtN4icUD4HCTt4B1Qmi3fj776GF8Qodghprag21x0bssdgIY3
AHDRU3PXoMaRcXXpCgNuqCSopJLzmzR/3nJvdNhrrqLvi9s+eGrupBfxfMlpilPO
+OZq165Yhdxq1xSTgYnYq08hXid71hQhEP4FpXcYXc7EQK1ZQggHYRSTEIuMh0rS
QlnzlswWHKewoQnRBIYT6x4UetoO488eev6yB+4eqJsgVMAYV2NjlYxyRgeZqg+p
RP/WmJTcuq7imDJJdVt73K4hrlr49DcXQv+atsHlDw6HSxeliPWHGDTQ7St4cScn
LAiKpYBjaL5O/dZ5r0lCel6d71Xtz0lKg//OH187GLbMhAOV+Kn0ZqTO2JmaWhuG
qMRWWFLGsYrFyV7h6adEuyLOTvJwKvvdkvsdnTtvUdEoNxVsGH1Yzdwzg7d/0uZZ
E4Vi1h3vkkGdxZ2QFtHtsYh6uL4nityBhm5cDtVI58kt2/6au1cjf6SLh2d7bgrT
2hdz7+mFVbMac70CQQ2sXUuyLY1QsriT0ixy7nrd1V8RU3IWVNIpViSVB6s/m0L2
FXqO79JruBRU3gVoJJD+dmtz+WWs7Wijz23voJpn4SSqPFcsuewykF2+BJOKLYNF
bMmC3gTX590E1AcAvoEDKdfQTz8RgtKFpLFvqwfoFy6TbXRKzc5QE9F7EgD1KFKr
MjrOcw1XOx284P7WB4YtJZVP9pkWlp8F4sroFz/WjGDbP2+Swr2UeXmSRQP2PjQp
ko3a2eLXIbA7RiFXFmRnpPF65SEfwOmiCqx/70i0n7/fFtgRYOCcWKEmtSY2wX39
UDxpWv1Odx9mi5PQZWGfAtxhcGcIrUtBQ6w0MNcwQwbq9OGghNVcwqZEl1ddvDTu
W7U0L+C8XztfYfGdQ8RMIJhlMjBkSGa3fhfIDGF+nrThBGF1UE9AcRAVcnYdnFyz
20CsCFflJ0tng+wW0Jrk+IzWIIvKgsK24tf3hYdy/JcqWSN3PZ4ofirF3POYqc4f
o9dPOGLK4KNFG1Ic3cyg7FQOO/pssnwe1QEYsRhZvyCMMqh45cPU0dxaqRffWNgD
QsfwRzWBUkx+Q8foAwxz/8JaNCNDMbIJko1Jp22nx7E=
//pragma protect end_data_block
//pragma protect digest_block
ozm2hedMr0i1GIRWPZzhmIJQZ7M=
//pragma protect end_digest_block
//pragma protect end_protected
