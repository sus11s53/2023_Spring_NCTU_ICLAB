//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
aWSuatfPMLAcd2Ur+e3fgKc8eZJ+dnYMcHgPe50rw0H5ImOlPMOnQX0caHc2xooL
2HCSf9vf0NxO6HKZtIFtziw4jiloVl2jdkbaCe6YOjDz0diU+qdOaJ8MedWRDg4Q
2qoYxh60GCj61LF6SZ/WX3IbrZLzaSVM6x7ocy9JMlbxufsXzAPYEbNRij7d1fI/
ILKbWCEph6zUdPlVTPN573H9ATKpGGPfxP0sU3H2oar0xo7DveBbThvqOB2ycAhJ
oCv15xxdfYat/1+HDRmIgf7gqzjQ4TksMSQycdQqjD4qudTlfEMpbsNsqHe7F8Ce
FUZytrOJgg4dzbT1iplD1Q==
//pragma protect end_key_block
//pragma protect digest_block
s6QsMDckJDlMl0Z9QPVVhiM7dSo=
//pragma protect end_digest_block
//pragma protect data_block
Gt5+MOx3+TP+HsCg677HfAlz360dugPYs0wEFSlu+DmuA1kPLYV6aVRQKf1DFZ+N
ZmuPVvXXI63slb4wJY6aUr8ezALezp0rEg4RmxzJFsUtbHrPcSOGW8MmjNsDi93T
fu5y3woJwEkiPCV8X8kwQN9DtP3jH9pns95Ikf9TKTNdUFAXvu8YK+XARH1ukrPA
THM3z4k/aTtfH0MGcBVhalxJ2rCtfxjC/2kCXN5efzi35R060KIn8oQxkZRT2yPS
0v1h1NyRw09umEyahk5mlOu4XfcHwYaZIQn20OYJ750upyayKEKvDKpbQ37P74JI
pZyyqVWNUTDIQ3S0XSLUufjEAs6y1ckQGhxaqmkKlwOUX53yxOblZqesdyKXdeK8
txW4wJPBcUmoUu6t6rpT0KFCESZVfvIjD/EH5oRjgf5BAEM4UnxzdOK8yh6Vh+o1
eUBaJ5XlVU7kNz9c5bFaDWro16uNZhQz1qI74ngZHSpyatwDIm4o5Hv0P1ceLh+b
co4FGDA1M8d2MtoCW7NRbvBNWzO/hklrBjkOzpH4JIuSHnK8hQ/hvx/WDT3imXk/
vLQ/8NIGjvkntUneQ6euft6abAeHAigmd4XCR7pC5INPH6mL4wlyNmgRKw3TeYdN
yfPSswRiaWf5nyXI1dWm9K3TG/smWJ1WKnko4uQGjWUq/pcEM0lu2FRM0gnb4x9f
nrLcmtwPeExLhsukqV3HteOa6KoLRdayqtM6HrBOshYZ4w4DjDIuYnjrjtoVZlNE
gYiGhzfRtBD+8mDvkC4W8wYWUAIW+C2iOZaML5Ya6mcFN2BuyjfWXaixg6zTxMq9
kQ1tbjZMCvFKYGmi+h3lr7yQODGDufcdZ8RwtATwtvHlcIfwx8U7WBKv1Wrwa/vx
QGUmO/peTubR455WwpiTYLeKkbHWGm9NhP8KLfmGxa3snS66MtZ9C4ICOQ7MufM8
tnhktKmqNUdxhZ2TH62PNpCS8rFkad/mh29eBNGiYGbJ3LKu2vYUJa/yvWGu+K59
7cemgIJnkwNFeXO7fxuutBJF14osI91lJIBfDh2O+2u/8oE17IzbZcyM8wime9hc
J6TZjbvw6J5xvRfv+K6jLqoVFdsvt19Bk/KUCmkkaK8sDPje9AShBT5wSyC5jDcu
sVsslq/1FDJ3PhFyh5XuvyfCliI6Xg6ZMhrOXsWYXoufh2vNmEM8zYG5ADPZVYS6
Taxovyq+AVwK4kOQYM7lAYGnEufLR5H+YEetZ+yykJsDRyG78vE/FW0GUy5QBh/C
ZyHahRPy6FK49q4PwUeuVFKAZmHAdaF4Lc7v+KmLJg6zNwQVtXunhvCt/Ityyxte
AOc/qVZUTMCHcUvaTGdK9K52sli5N6mk52x6G1zXSHmVF3N3VQVkEok2AyTQRl25
t7TMPrZ+VxW5eX/h49bShBWQ7sR1JWcuOLPYsQtYfBDDVPPrEh5DGL/z6rGcpzfk
KUjTy0k2ftlq4yLS74SNar9AqZ5odKM6iD+C9v7E5rjV/SG+7q0CkaFBUp5zuwdc
cmD4LeFQMx2r+d/pWdLtH4eBdZ1earVwkrk+KUND6TnjBFhxYRBwkC9xGALnb6n4
pWRqmDre9FeqBho0Kh3gup3n1n/m/bAEq3QyGPO+McIOaOzeTtq+I0NizokaZ5/V
NwR0ji4VtndWMXNDj2aMbVyMeOzRVObcNQOaPzbQGTH1S/ZyJNqYI/CHWoYzGn/u
XZSVrpV2P6TRWqu8IhSuKbLXil2MnOUnlDtp/SXHrezkVW1NJ1BAUbe8sRQuA3A5
kGECjMr0/VYQoUY4QsN54H2qGdaHDfG0433tp7ryYzB/kNeP1bhKHxbQ9RLX7gdK
qZgB6NtNdvabSwaUvTRfDEde7abSvUa80u5RfMlqhHLGHtAo+id0eQHOoCZwLJwM
SjI+kVk4opYK8P3jIm5AJ6doxmrfTD3C3uLCFbTYt6T0YwDPy6IdGH55+ukt0iKd
IZUYmnyQAmNb60WM8DfUm9poRuHMvhENuL3+VvsBuQDQiIPn9WmSsDhaniWYm1Yq
5toe0r+gS6o8X3AnL2cPznOZ1IDWCSfA02Lz87LKUJJOmclAQ7lKdOVSD4TxWf/o
4D9WPigGTnruGNoqFOWOoH958f9B6ILPspTuWztl0KplsxOwHuNGY9qDnPEMVZxI
wBM17gz0xfc8iWLUllLbLb6PB98pQIwXyyfcJnti1VoBFtk4xPt8u1NOtzZyK4vR
u2mxQ5nuTrHPcKCTGlP0SibeuBismo9c1JlxfLh1XRbs8/ZcXGGJMjX1MjZ6BH/k
7KijoW1uEvHf87zEQjIM3Di44KlrhBPOu8E37DpBUb3tNEuTvye+AboHDn2LEFDz
6drDx248172/kkFGRjpPHdpj9Z0QN9U0n0oXSP4OxF2SHhaAP0TuRYi+kYtSp+nn
rp4M38iHu6fn6K504dmecgchZ+qZwAshbT5GqR509XNCkY6dSyaYceMD4WxXlqzy
PE03Ym6vHyiBUmpTP8HKgR0OmZ/LqqV5mlKdwI7iVUhvZSiz4A90DjyvFXP1rwtH
Wd3smTppJKW7VxB1V9jbCd+MGp9EnNqgVSOP9NE0upQefZ7RcLNP8W71BfhmAeUa
EnJtF9JBTICSQqpbIv/sajUBh45aLvvgQf+fBZxn8aWTF9uKTVbopfIQRjj+rGVZ
03iWGLTm8fSgmb3HahKFGhWIjmuoT5m1uOd+tiwsPLeqMUEm+NNZbniSE0vTPT91
yUe9lCm/FAXlaCl6egcDbFtBIdBuHFZOyqP7a2UI/oFS8yd6gcCfXpCq0b/EzKo6
lzStoBKZhphxRnW4rBJ5PsgBJw/toeZOr0PiBUheIoS8/Uz4/19rwwHx7nPhFKnW
9INoD5jiAeUXareUGUOij7ktDWW0Gb/qKhVlUly4WZA3PzGzZoQjZ3P7znJxrNBy
oQDKZ7+xEDErhqrsJM6rjyh7+hnsNbg4Ndy4d1zR05E8mlFt1OrwunA+es4BR/7U
71/LPy7JwrSTGNY+zBAZ5RUbDSynnzQwZBEbHpsgRwla1MB9GpvlXfiS22jAScTo
QKLKwhv7gpi5d600LDtc4plplYweVOqsZu6arh9P+amQ1yRqFujnos60ygOZz1gn
uxu94c1kVfpgQd1rNSMLUJyGOZwdDeRbbujnqsTdztfFw0fFUthRRKcDay37sIGV
dQz6qkKjouWhA12FWOAADhBATb3evg69UlddhTwVBGjtLyUthXa6WkWGmzkMb5lo
zHVdckPz+NfKnBQAC7sx/U7SD9+2IzyMm6G6vH8MQuNh5egLuDQx0dkpp4CqXove
7L9+0ctpgmoRwtsLswWHlGP3dgBE1kM48svO24I2/+QA6KyH4UhMpVN6BZ4bSKwN
jkP67GiZq+oPRe36cuQAFHxfAzYAmkCtD5KiuAZz1SVOQHe4Y4nV8YGNIKZ5sTxx
od1L51Nkyb0sls+pKsDI+EUukX0mUHsiGs8HncRjH84=
//pragma protect end_data_block
//pragma protect digest_block
TufOJhiv+TCQCSI8R7u5Omj5Bo8=
//pragma protect end_digest_block
//pragma protect end_protected
